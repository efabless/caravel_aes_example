VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aes_example
  CLASS BLOCK ;
  FOREIGN aes_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 820.000 BY 800.000 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 795.440 10.640 798.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 713.840 10.640 717.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.240 10.640 635.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.640 10.640 553.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.040 10.640 472.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.440 10.640 390.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 305.840 10.640 309.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.240 10.640 227.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 142.640 10.640 145.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.040 10.640 64.240 789.040 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 754.640 10.640 757.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 673.040 10.640 676.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.440 10.640 594.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 509.840 10.640 513.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.240 10.640 431.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.640 10.640 349.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 265.040 10.640 268.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.440 10.640 186.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.840 10.640 105.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.240 10.640 23.440 789.040 ;
    END
  END VPWR
  PIN wb_clk_i
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 751.730 0.000 752.010 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 784.665 814.390 787.495 ;
        RECT 5.330 779.225 814.390 782.055 ;
        RECT 5.330 773.785 814.390 776.615 ;
        RECT 5.330 768.345 814.390 771.175 ;
        RECT 5.330 762.905 814.390 765.735 ;
        RECT 5.330 757.465 814.390 760.295 ;
        RECT 5.330 752.025 814.390 754.855 ;
        RECT 5.330 746.585 814.390 749.415 ;
        RECT 5.330 741.145 814.390 743.975 ;
        RECT 5.330 735.705 814.390 738.535 ;
        RECT 5.330 730.265 814.390 733.095 ;
        RECT 5.330 724.825 814.390 727.655 ;
        RECT 5.330 719.385 814.390 722.215 ;
        RECT 5.330 713.945 814.390 716.775 ;
        RECT 5.330 708.505 814.390 711.335 ;
        RECT 5.330 703.065 814.390 705.895 ;
        RECT 5.330 697.625 814.390 700.455 ;
        RECT 5.330 692.185 814.390 695.015 ;
        RECT 5.330 686.745 814.390 689.575 ;
        RECT 5.330 681.305 814.390 684.135 ;
        RECT 5.330 675.865 814.390 678.695 ;
        RECT 5.330 670.425 814.390 673.255 ;
        RECT 5.330 664.985 814.390 667.815 ;
        RECT 5.330 659.545 814.390 662.375 ;
        RECT 5.330 654.105 814.390 656.935 ;
        RECT 5.330 648.665 814.390 651.495 ;
        RECT 5.330 643.225 814.390 646.055 ;
        RECT 5.330 637.785 814.390 640.615 ;
        RECT 5.330 632.345 814.390 635.175 ;
        RECT 5.330 626.905 814.390 629.735 ;
        RECT 5.330 621.465 814.390 624.295 ;
        RECT 5.330 616.025 814.390 618.855 ;
        RECT 5.330 610.585 814.390 613.415 ;
        RECT 5.330 605.145 814.390 607.975 ;
        RECT 5.330 599.705 814.390 602.535 ;
        RECT 5.330 594.265 814.390 597.095 ;
        RECT 5.330 588.825 814.390 591.655 ;
        RECT 5.330 583.385 814.390 586.215 ;
        RECT 5.330 577.945 814.390 580.775 ;
        RECT 5.330 572.505 814.390 575.335 ;
        RECT 5.330 567.065 814.390 569.895 ;
        RECT 5.330 561.625 814.390 564.455 ;
        RECT 5.330 556.185 814.390 559.015 ;
        RECT 5.330 550.745 814.390 553.575 ;
        RECT 5.330 545.305 814.390 548.135 ;
        RECT 5.330 539.865 814.390 542.695 ;
        RECT 5.330 534.425 814.390 537.255 ;
        RECT 5.330 528.985 814.390 531.815 ;
        RECT 5.330 523.545 814.390 526.375 ;
        RECT 5.330 518.105 814.390 520.935 ;
        RECT 5.330 512.665 814.390 515.495 ;
        RECT 5.330 507.225 814.390 510.055 ;
        RECT 5.330 501.785 814.390 504.615 ;
        RECT 5.330 496.345 814.390 499.175 ;
        RECT 5.330 490.905 814.390 493.735 ;
        RECT 5.330 485.465 814.390 488.295 ;
        RECT 5.330 480.025 814.390 482.855 ;
        RECT 5.330 474.585 814.390 477.415 ;
        RECT 5.330 469.145 814.390 471.975 ;
        RECT 5.330 463.705 814.390 466.535 ;
        RECT 5.330 458.265 814.390 461.095 ;
        RECT 5.330 452.825 814.390 455.655 ;
        RECT 5.330 447.385 814.390 450.215 ;
        RECT 5.330 441.945 814.390 444.775 ;
        RECT 5.330 436.505 814.390 439.335 ;
        RECT 5.330 431.065 814.390 433.895 ;
        RECT 5.330 425.625 814.390 428.455 ;
        RECT 5.330 420.185 814.390 423.015 ;
        RECT 5.330 414.745 814.390 417.575 ;
        RECT 5.330 409.305 814.390 412.135 ;
        RECT 5.330 403.865 814.390 406.695 ;
        RECT 5.330 398.425 814.390 401.255 ;
        RECT 5.330 392.985 814.390 395.815 ;
        RECT 5.330 387.545 814.390 390.375 ;
        RECT 5.330 382.105 814.390 384.935 ;
        RECT 5.330 376.665 814.390 379.495 ;
        RECT 5.330 371.225 814.390 374.055 ;
        RECT 5.330 365.785 814.390 368.615 ;
        RECT 5.330 360.345 814.390 363.175 ;
        RECT 5.330 354.905 814.390 357.735 ;
        RECT 5.330 349.465 814.390 352.295 ;
        RECT 5.330 344.025 814.390 346.855 ;
        RECT 5.330 338.585 814.390 341.415 ;
        RECT 5.330 333.145 814.390 335.975 ;
        RECT 5.330 327.705 814.390 330.535 ;
        RECT 5.330 322.265 814.390 325.095 ;
        RECT 5.330 316.825 814.390 319.655 ;
        RECT 5.330 311.385 814.390 314.215 ;
        RECT 5.330 305.945 814.390 308.775 ;
        RECT 5.330 300.505 814.390 303.335 ;
        RECT 5.330 295.065 814.390 297.895 ;
        RECT 5.330 289.625 814.390 292.455 ;
        RECT 5.330 284.185 814.390 287.015 ;
        RECT 5.330 278.745 814.390 281.575 ;
        RECT 5.330 273.305 814.390 276.135 ;
        RECT 5.330 267.865 814.390 270.695 ;
        RECT 5.330 262.425 814.390 265.255 ;
        RECT 5.330 256.985 814.390 259.815 ;
        RECT 5.330 251.545 814.390 254.375 ;
        RECT 5.330 246.105 814.390 248.935 ;
        RECT 5.330 240.665 814.390 243.495 ;
        RECT 5.330 235.225 814.390 238.055 ;
        RECT 5.330 229.785 814.390 232.615 ;
        RECT 5.330 224.345 814.390 227.175 ;
        RECT 5.330 218.905 814.390 221.735 ;
        RECT 5.330 213.465 814.390 216.295 ;
        RECT 5.330 208.025 814.390 210.855 ;
        RECT 5.330 202.585 814.390 205.415 ;
        RECT 5.330 197.145 814.390 199.975 ;
        RECT 5.330 191.705 814.390 194.535 ;
        RECT 5.330 186.265 814.390 189.095 ;
        RECT 5.330 180.825 814.390 183.655 ;
        RECT 5.330 175.385 814.390 178.215 ;
        RECT 5.330 169.945 814.390 172.775 ;
        RECT 5.330 164.505 814.390 167.335 ;
        RECT 5.330 159.065 814.390 161.895 ;
        RECT 5.330 153.625 814.390 156.455 ;
        RECT 5.330 148.185 814.390 151.015 ;
        RECT 5.330 142.745 814.390 145.575 ;
        RECT 5.330 137.305 814.390 140.135 ;
        RECT 5.330 131.865 814.390 134.695 ;
        RECT 5.330 126.425 814.390 129.255 ;
        RECT 5.330 120.985 814.390 123.815 ;
        RECT 5.330 115.545 814.390 118.375 ;
        RECT 5.330 110.105 814.390 112.935 ;
        RECT 5.330 104.665 814.390 107.495 ;
        RECT 5.330 99.225 814.390 102.055 ;
        RECT 5.330 93.785 814.390 96.615 ;
        RECT 5.330 88.345 814.390 91.175 ;
        RECT 5.330 82.905 814.390 85.735 ;
        RECT 5.330 77.465 814.390 80.295 ;
        RECT 5.330 72.025 814.390 74.855 ;
        RECT 5.330 66.585 814.390 69.415 ;
        RECT 5.330 61.145 814.390 63.975 ;
        RECT 5.330 55.705 814.390 58.535 ;
        RECT 5.330 50.265 814.390 53.095 ;
        RECT 5.330 44.825 814.390 47.655 ;
        RECT 5.330 39.385 814.390 42.215 ;
        RECT 5.330 33.945 814.390 36.775 ;
        RECT 5.330 28.505 814.390 31.335 ;
        RECT 5.330 23.065 814.390 25.895 ;
        RECT 5.330 17.625 814.390 20.455 ;
        RECT 5.330 12.185 814.390 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 814.200 788.885 ;
      LAYER met1 ;
        RECT 5.520 4.120 815.050 789.040 ;
      LAYER met2 ;
        RECT 7.000 4.280 815.020 788.985 ;
        RECT 7.000 3.555 22.810 4.280 ;
        RECT 23.650 3.555 30.170 4.280 ;
        RECT 31.010 3.555 37.530 4.280 ;
        RECT 38.370 3.555 44.890 4.280 ;
        RECT 45.730 3.555 52.250 4.280 ;
        RECT 53.090 3.555 59.610 4.280 ;
        RECT 60.450 3.555 66.970 4.280 ;
        RECT 67.810 3.555 74.330 4.280 ;
        RECT 75.170 3.555 81.690 4.280 ;
        RECT 82.530 3.555 89.050 4.280 ;
        RECT 89.890 3.555 96.410 4.280 ;
        RECT 97.250 3.555 103.770 4.280 ;
        RECT 104.610 3.555 111.130 4.280 ;
        RECT 111.970 3.555 118.490 4.280 ;
        RECT 119.330 3.555 125.850 4.280 ;
        RECT 126.690 3.555 133.210 4.280 ;
        RECT 134.050 3.555 140.570 4.280 ;
        RECT 141.410 3.555 147.930 4.280 ;
        RECT 148.770 3.555 155.290 4.280 ;
        RECT 156.130 3.555 162.650 4.280 ;
        RECT 163.490 3.555 170.010 4.280 ;
        RECT 170.850 3.555 177.370 4.280 ;
        RECT 178.210 3.555 184.730 4.280 ;
        RECT 185.570 3.555 192.090 4.280 ;
        RECT 192.930 3.555 199.450 4.280 ;
        RECT 200.290 3.555 206.810 4.280 ;
        RECT 207.650 3.555 214.170 4.280 ;
        RECT 215.010 3.555 221.530 4.280 ;
        RECT 222.370 3.555 228.890 4.280 ;
        RECT 229.730 3.555 236.250 4.280 ;
        RECT 237.090 3.555 243.610 4.280 ;
        RECT 244.450 3.555 250.970 4.280 ;
        RECT 251.810 3.555 258.330 4.280 ;
        RECT 259.170 3.555 265.690 4.280 ;
        RECT 266.530 3.555 273.050 4.280 ;
        RECT 273.890 3.555 280.410 4.280 ;
        RECT 281.250 3.555 287.770 4.280 ;
        RECT 288.610 3.555 295.130 4.280 ;
        RECT 295.970 3.555 302.490 4.280 ;
        RECT 303.330 3.555 309.850 4.280 ;
        RECT 310.690 3.555 317.210 4.280 ;
        RECT 318.050 3.555 324.570 4.280 ;
        RECT 325.410 3.555 331.930 4.280 ;
        RECT 332.770 3.555 339.290 4.280 ;
        RECT 340.130 3.555 346.650 4.280 ;
        RECT 347.490 3.555 354.010 4.280 ;
        RECT 354.850 3.555 361.370 4.280 ;
        RECT 362.210 3.555 368.730 4.280 ;
        RECT 369.570 3.555 376.090 4.280 ;
        RECT 376.930 3.555 383.450 4.280 ;
        RECT 384.290 3.555 390.810 4.280 ;
        RECT 391.650 3.555 398.170 4.280 ;
        RECT 399.010 3.555 405.530 4.280 ;
        RECT 406.370 3.555 412.890 4.280 ;
        RECT 413.730 3.555 420.250 4.280 ;
        RECT 421.090 3.555 427.610 4.280 ;
        RECT 428.450 3.555 434.970 4.280 ;
        RECT 435.810 3.555 442.330 4.280 ;
        RECT 443.170 3.555 449.690 4.280 ;
        RECT 450.530 3.555 457.050 4.280 ;
        RECT 457.890 3.555 464.410 4.280 ;
        RECT 465.250 3.555 471.770 4.280 ;
        RECT 472.610 3.555 479.130 4.280 ;
        RECT 479.970 3.555 486.490 4.280 ;
        RECT 487.330 3.555 493.850 4.280 ;
        RECT 494.690 3.555 501.210 4.280 ;
        RECT 502.050 3.555 508.570 4.280 ;
        RECT 509.410 3.555 515.930 4.280 ;
        RECT 516.770 3.555 523.290 4.280 ;
        RECT 524.130 3.555 530.650 4.280 ;
        RECT 531.490 3.555 538.010 4.280 ;
        RECT 538.850 3.555 545.370 4.280 ;
        RECT 546.210 3.555 552.730 4.280 ;
        RECT 553.570 3.555 560.090 4.280 ;
        RECT 560.930 3.555 567.450 4.280 ;
        RECT 568.290 3.555 574.810 4.280 ;
        RECT 575.650 3.555 582.170 4.280 ;
        RECT 583.010 3.555 589.530 4.280 ;
        RECT 590.370 3.555 596.890 4.280 ;
        RECT 597.730 3.555 604.250 4.280 ;
        RECT 605.090 3.555 611.610 4.280 ;
        RECT 612.450 3.555 618.970 4.280 ;
        RECT 619.810 3.555 626.330 4.280 ;
        RECT 627.170 3.555 633.690 4.280 ;
        RECT 634.530 3.555 641.050 4.280 ;
        RECT 641.890 3.555 648.410 4.280 ;
        RECT 649.250 3.555 655.770 4.280 ;
        RECT 656.610 3.555 663.130 4.280 ;
        RECT 663.970 3.555 670.490 4.280 ;
        RECT 671.330 3.555 677.850 4.280 ;
        RECT 678.690 3.555 685.210 4.280 ;
        RECT 686.050 3.555 692.570 4.280 ;
        RECT 693.410 3.555 699.930 4.280 ;
        RECT 700.770 3.555 707.290 4.280 ;
        RECT 708.130 3.555 714.650 4.280 ;
        RECT 715.490 3.555 722.010 4.280 ;
        RECT 722.850 3.555 729.370 4.280 ;
        RECT 730.210 3.555 736.730 4.280 ;
        RECT 737.570 3.555 744.090 4.280 ;
        RECT 744.930 3.555 751.450 4.280 ;
        RECT 752.290 3.555 758.810 4.280 ;
        RECT 759.650 3.555 766.170 4.280 ;
        RECT 767.010 3.555 773.530 4.280 ;
        RECT 774.370 3.555 780.890 4.280 ;
        RECT 781.730 3.555 788.250 4.280 ;
        RECT 789.090 3.555 795.610 4.280 ;
        RECT 796.450 3.555 815.020 4.280 ;
      LAYER met3 ;
        RECT 19.845 3.575 813.215 788.965 ;
      LAYER met4 ;
        RECT 30.655 10.240 60.640 735.585 ;
        RECT 64.640 10.240 101.440 735.585 ;
        RECT 105.440 10.240 142.240 735.585 ;
        RECT 146.240 10.240 183.040 735.585 ;
        RECT 187.040 10.240 223.840 735.585 ;
        RECT 227.840 10.240 264.640 735.585 ;
        RECT 268.640 10.240 305.440 735.585 ;
        RECT 309.440 10.240 346.240 735.585 ;
        RECT 350.240 10.240 387.040 735.585 ;
        RECT 391.040 10.240 427.840 735.585 ;
        RECT 431.840 10.240 468.640 735.585 ;
        RECT 472.640 10.240 509.440 735.585 ;
        RECT 513.440 10.240 550.240 735.585 ;
        RECT 554.240 10.240 591.040 735.585 ;
        RECT 595.040 10.240 631.840 735.585 ;
        RECT 635.840 10.240 672.640 735.585 ;
        RECT 676.640 10.240 713.440 735.585 ;
        RECT 717.440 10.240 754.240 735.585 ;
        RECT 758.240 10.240 795.040 735.585 ;
        RECT 799.040 10.240 804.705 735.585 ;
        RECT 30.655 3.575 804.705 10.240 ;
  END
END aes_example
END LIBRARY

