magic
tech sky130A
magscale 1 2
timestamp 1686002167
<< obsli1 >>
rect 3104 6159 164840 161777
<< obsm1 >>
rect 3104 2048 165010 161808
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 570 536 165004 161797
rect 710 326 1590 536
rect 1814 326 2786 536
rect 3010 326 3982 536
rect 4206 326 5178 536
rect 5402 326 6374 536
rect 6598 326 7570 536
rect 7794 326 8674 536
rect 8898 326 9870 536
rect 10094 326 11066 536
rect 11290 326 12262 536
rect 12486 326 13458 536
rect 13682 326 14654 536
rect 14878 326 15850 536
rect 16074 326 16954 536
rect 17178 326 18150 536
rect 18374 326 19346 536
rect 19570 326 20542 536
rect 20766 326 21738 536
rect 21962 326 22934 536
rect 23158 326 24130 536
rect 24354 326 25234 536
rect 25458 326 26430 536
rect 26654 326 27626 536
rect 27850 326 28822 536
rect 29046 326 30018 536
rect 30242 326 31214 536
rect 31438 326 32318 536
rect 32542 326 33514 536
rect 33738 326 34710 536
rect 34934 326 35906 536
rect 36130 326 37102 536
rect 37326 326 38298 536
rect 38522 326 39494 536
rect 39718 326 40598 536
rect 40822 326 41794 536
rect 42018 326 42990 536
rect 43214 326 44186 536
rect 44410 326 45382 536
rect 45606 326 46578 536
rect 46802 326 47774 536
rect 47998 326 48878 536
rect 49102 326 50074 536
rect 50298 326 51270 536
rect 51494 326 52466 536
rect 52690 326 53662 536
rect 53886 326 54858 536
rect 55082 326 55962 536
rect 56186 326 57158 536
rect 57382 326 58354 536
rect 58578 326 59550 536
rect 59774 326 60746 536
rect 60970 326 61942 536
rect 62166 326 63138 536
rect 63362 326 64242 536
rect 64466 326 65438 536
rect 65662 326 66634 536
rect 66858 326 67830 536
rect 68054 326 69026 536
rect 69250 326 70222 536
rect 70446 326 71418 536
rect 71642 326 72522 536
rect 72746 326 73718 536
rect 73942 326 74914 536
rect 75138 326 76110 536
rect 76334 326 77306 536
rect 77530 326 78502 536
rect 78726 326 79606 536
rect 79830 326 80802 536
rect 81026 326 81998 536
rect 82222 326 83194 536
rect 83418 326 84390 536
rect 84614 326 85586 536
rect 85810 326 86782 536
rect 87006 326 87886 536
rect 88110 326 89082 536
rect 89306 326 90278 536
rect 90502 326 91474 536
rect 91698 326 92670 536
rect 92894 326 93866 536
rect 94090 326 95062 536
rect 95286 326 96166 536
rect 96390 326 97362 536
rect 97586 326 98558 536
rect 98782 326 99754 536
rect 99978 326 100950 536
rect 101174 326 102146 536
rect 102370 326 103250 536
rect 103474 326 104446 536
rect 104670 326 105642 536
rect 105866 326 106838 536
rect 107062 326 108034 536
rect 108258 326 109230 536
rect 109454 326 110426 536
rect 110650 326 111530 536
rect 111754 326 112726 536
rect 112950 326 113922 536
rect 114146 326 115118 536
rect 115342 326 116314 536
rect 116538 326 117510 536
rect 117734 326 118706 536
rect 118930 326 119810 536
rect 120034 326 121006 536
rect 121230 326 122202 536
rect 122426 326 123398 536
rect 123622 326 124594 536
rect 124818 326 125790 536
rect 126014 326 126894 536
rect 127118 326 128090 536
rect 128314 326 129286 536
rect 129510 326 130482 536
rect 130706 326 131678 536
rect 131902 326 132874 536
rect 133098 326 134070 536
rect 134294 326 135174 536
rect 135398 326 136370 536
rect 136594 326 137566 536
rect 137790 326 138762 536
rect 138986 326 139958 536
rect 140182 326 141154 536
rect 141378 326 142350 536
rect 142574 326 143454 536
rect 143678 326 144650 536
rect 144874 326 145846 536
rect 146070 326 147042 536
rect 147266 326 148238 536
rect 148462 326 149434 536
rect 149658 326 150538 536
rect 150762 326 151734 536
rect 151958 326 152930 536
rect 153154 326 154126 536
rect 154350 326 155322 536
rect 155546 326 156518 536
rect 156742 326 157714 536
rect 157938 326 158818 536
rect 159042 326 160014 536
rect 160238 326 161210 536
rect 161434 326 162406 536
rect 162630 326 163602 536
rect 163826 326 164798 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect -960 149684 480 149924
rect -960 136628 480 136868
rect -960 123572 480 123812
rect -960 110516 480 110756
rect -960 97460 480 97700
rect -960 84540 480 84780
rect -960 71484 480 71724
rect -960 58428 480 58668
rect -960 45372 480 45612
rect -960 32316 480 32556
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 152540 584960 152780
rect 583520 139212 584960 139452
rect 583520 125884 584960 126124
rect 583520 112692 584960 112932
rect 583520 99364 584960 99604
rect 583520 86036 584960 86276
rect 583520 72844 584960 73084
rect 583520 59516 584960 59756
rect 583520 46188 584960 46428
rect 583520 32996 584960 33236
rect 583520 19668 584960 19908
rect 583520 6476 584960 6716
<< obsm3 >>
rect 565 1667 164643 161793
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1784 -7654 2424 711590
rect 3064 -7654 3704 711590
rect 4344 -7654 4984 711590
rect 5624 161888 6264 711590
rect 6904 151257 7544 711590
rect 8184 151257 8824 711590
rect 9464 151257 10104 711590
rect 10744 151257 11384 711590
rect 18104 151257 18744 711590
rect 19384 151257 20024 711590
rect 20664 151257 21304 711590
rect 21944 161888 22584 711590
rect 23224 151257 23864 711590
rect 24504 151257 25144 711590
rect 25784 151257 26424 711590
rect 27064 151257 27704 711590
rect 34424 151257 35064 711590
rect 35704 151257 36344 711590
rect 36984 151257 37624 711590
rect 38264 161888 38904 711590
rect 39544 151257 40184 711590
rect 40824 151257 41464 711590
rect 42104 151257 42744 711590
rect 43384 151257 44024 711590
rect 50744 151257 51384 711590
rect 52024 151257 52664 711590
rect 53304 151257 53944 711590
rect 54584 161888 55224 711590
rect 55864 151257 56504 711590
rect 57144 151257 57784 711590
rect 58424 151257 59064 711590
rect 59704 151257 60344 711590
rect 67064 151257 67704 711590
rect 68344 151257 68984 711590
rect 69624 151257 70264 711590
rect 70904 161888 71544 711590
rect 72184 151257 72824 711590
rect 73464 151257 74104 711590
rect 74744 151257 75384 711590
rect 76024 151257 76664 711590
rect 83384 151257 84024 711590
rect 84664 151257 85304 711590
rect 85944 151257 86584 711590
rect 87224 161888 87864 711590
rect 88504 151257 89144 711590
rect 89784 151257 90424 711590
rect 91064 151257 91704 711590
rect 92344 151257 92984 711590
rect 99704 151257 100344 711590
rect 100984 151257 101624 711590
rect 102264 151257 102904 711590
rect 103544 161888 104184 711590
rect 104824 151257 105464 711590
rect 106104 151257 106744 711590
rect 107384 151257 108024 711590
rect 108664 151257 109304 711590
rect 116024 151257 116664 711590
rect 117304 151257 117944 711590
rect 118584 151257 119224 711590
rect 119864 161888 120504 711590
rect 121144 151257 121784 711590
rect 122424 151257 123064 711590
rect 123704 151257 124344 711590
rect 124984 151257 125624 711590
rect 132344 151257 132984 711590
rect 133624 151257 134264 711590
rect 134904 151257 135544 711590
rect 136184 161888 136824 711590
rect 137464 151257 138104 711590
rect 138744 151257 139384 711590
rect 140024 151257 140664 711590
rect 141304 151257 141944 711590
rect 148664 151257 149304 711590
rect 149944 151257 150584 711590
rect 151224 151257 151864 711590
rect 152504 161888 153144 711590
rect 153784 151257 154424 711590
rect 155064 151257 155704 711590
rect 156344 151257 156984 711590
rect 157624 151257 158264 711590
rect 164984 151257 165624 711590
rect 18104 -7654 18744 4575
rect 19384 -7654 20024 4575
rect 34424 -7654 35064 4575
rect 35704 -7654 36344 4575
rect 50744 -7654 51384 4575
rect 52024 -7654 52664 4575
rect 67064 -7654 67704 4575
rect 68344 -7654 68984 4575
rect 83384 -7654 84024 4575
rect 84664 -7654 85304 4575
rect 99704 -7654 100344 4575
rect 100984 -7654 101624 4575
rect 116024 -7654 116664 4575
rect 117304 -7654 117944 4575
rect 132344 -7654 132984 4575
rect 133624 -7654 134264 4575
rect 148664 -7654 149304 4575
rect 149944 -7654 150584 4575
rect 164984 -7654 165624 4575
rect 166264 -7654 166904 711590
rect 167544 -7654 168184 711590
rect 168824 -7654 169464 711590
rect 170104 -7654 170744 711590
rect 171384 -7654 172024 711590
rect 172664 -7654 173304 711590
rect 173944 -7654 174584 711590
rect 181304 -7654 181944 711590
rect 182584 -7654 183224 711590
rect 183864 -7654 184504 711590
rect 185144 -7654 185784 711590
rect 186424 -7654 187064 711590
rect 187704 -7654 188344 711590
rect 188984 -7654 189624 711590
rect 190264 -7654 190904 711590
rect 197624 -7654 198264 711590
rect 198904 -7654 199544 711590
rect 200184 -7654 200824 711590
rect 201464 -7654 202104 711590
rect 202744 -7654 203384 711590
rect 204024 -7654 204664 711590
rect 205304 -7654 205944 711590
rect 206584 -7654 207224 711590
rect 213944 -7654 214584 711590
rect 215224 -7654 215864 711590
rect 216504 -7654 217144 711590
rect 217784 -7654 218424 711590
rect 219064 -7654 219704 711590
rect 220344 -7654 220984 711590
rect 221624 -7654 222264 711590
rect 222904 -7654 223544 711590
rect 230264 -7654 230904 711590
rect 231544 -7654 232184 711590
rect 232824 -7654 233464 711590
rect 234104 -7654 234744 711590
rect 235384 -7654 236024 711590
rect 236664 -7654 237304 711590
rect 237944 -7654 238584 711590
rect 239224 -7654 239864 711590
rect 246584 -7654 247224 711590
rect 247864 -7654 248504 711590
rect 249144 -7654 249784 711590
rect 250424 -7654 251064 711590
rect 251704 -7654 252344 711590
rect 252984 -7654 253624 711590
rect 254264 -7654 254904 711590
rect 255544 -7654 256184 711590
rect 262904 -7654 263544 711590
rect 264184 -7654 264824 711590
rect 265464 -7654 266104 711590
rect 266744 -7654 267384 711590
rect 268024 -7654 268664 711590
rect 269304 -7654 269944 711590
rect 270584 -7654 271224 711590
rect 271864 -7654 272504 711590
rect 279224 -7654 279864 711590
rect 280504 -7654 281144 711590
rect 281784 -7654 282424 711590
rect 283064 -7654 283704 711590
rect 284344 -7654 284984 711590
rect 285624 -7654 286264 711590
rect 286904 -7654 287544 711590
rect 288184 -7654 288824 711590
rect 295544 -7654 296184 711590
rect 296824 -7654 297464 711590
rect 298104 -7654 298744 711590
rect 299384 -7654 300024 711590
rect 300664 -7654 301304 711590
rect 301944 -7654 302584 711590
rect 303224 -7654 303864 711590
rect 304504 -7654 305144 711590
rect 311864 -7654 312504 711590
rect 313144 -7654 313784 711590
rect 314424 -7654 315064 711590
rect 315704 -7654 316344 711590
rect 316984 -7654 317624 711590
rect 318264 -7654 318904 711590
rect 319544 -7654 320184 711590
rect 320824 -7654 321464 711590
rect 328184 -7654 328824 711590
rect 329464 -7654 330104 711590
rect 330744 -7654 331384 711590
rect 332024 -7654 332664 711590
rect 333304 -7654 333944 711590
rect 334584 -7654 335224 711590
rect 335864 -7654 336504 711590
rect 337144 -7654 337784 711590
rect 344504 -7654 345144 711590
rect 345784 -7654 346424 711590
rect 347064 -7654 347704 711590
rect 348344 -7654 348984 711590
rect 349624 -7654 350264 711590
rect 350904 -7654 351544 711590
rect 352184 -7654 352824 711590
rect 353464 -7654 354104 711590
rect 360824 -7654 361464 711590
rect 362104 -7654 362744 711590
rect 363384 -7654 364024 711590
rect 364664 -7654 365304 711590
rect 365944 -7654 366584 711590
rect 367224 -7654 367864 711590
rect 368504 -7654 369144 711590
rect 369784 -7654 370424 711590
rect 377144 -7654 377784 711590
rect 378424 -7654 379064 711590
rect 379704 -7654 380344 711590
rect 380984 -7654 381624 711590
rect 382264 -7654 382904 711590
rect 383544 -7654 384184 711590
rect 384824 -7654 385464 711590
rect 386104 -7654 386744 711590
rect 393464 -7654 394104 711590
rect 394744 -7654 395384 711590
rect 396024 -7654 396664 711590
rect 397304 -7654 397944 711590
rect 398584 -7654 399224 711590
rect 399864 -7654 400504 711590
rect 401144 -7654 401784 711590
rect 402424 -7654 403064 711590
rect 409784 -7654 410424 711590
rect 411064 -7654 411704 711590
rect 412344 -7654 412984 711590
rect 413624 -7654 414264 711590
rect 414904 -7654 415544 711590
rect 416184 -7654 416824 711590
rect 417464 -7654 418104 711590
rect 418744 -7654 419384 711590
rect 426104 -7654 426744 711590
rect 427384 -7654 428024 711590
rect 428664 -7654 429304 711590
rect 429944 -7654 430584 711590
rect 431224 -7654 431864 711590
rect 432504 -7654 433144 711590
rect 433784 -7654 434424 711590
rect 435064 -7654 435704 711590
rect 442424 -7654 443064 711590
rect 443704 -7654 444344 711590
rect 444984 -7654 445624 711590
rect 446264 -7654 446904 711590
rect 447544 -7654 448184 711590
rect 448824 -7654 449464 711590
rect 450104 -7654 450744 711590
rect 451384 -7654 452024 711590
rect 458744 -7654 459384 711590
rect 460024 -7654 460664 711590
rect 461304 -7654 461944 711590
rect 462584 -7654 463224 711590
rect 463864 -7654 464504 711590
rect 465144 -7654 465784 711590
rect 466424 -7654 467064 711590
rect 467704 -7654 468344 711590
rect 475064 -7654 475704 711590
rect 476344 -7654 476984 711590
rect 477624 -7654 478264 711590
rect 478904 -7654 479544 711590
rect 480184 -7654 480824 711590
rect 481464 -7654 482104 711590
rect 482744 -7654 483384 711590
rect 484024 -7654 484664 711590
rect 491384 -7654 492024 711590
rect 492664 -7654 493304 711590
rect 493944 -7654 494584 711590
rect 495224 -7654 495864 711590
rect 496504 -7654 497144 711590
rect 497784 -7654 498424 711590
rect 499064 -7654 499704 711590
rect 500344 -7654 500984 711590
rect 507704 -7654 508344 711590
rect 508984 -7654 509624 711590
rect 510264 -7654 510904 711590
rect 511544 -7654 512184 711590
rect 512824 -7654 513464 711590
rect 514104 -7654 514744 711590
rect 515384 -7654 516024 711590
rect 516664 -7654 517304 711590
rect 524024 -7654 524664 711590
rect 525304 -7654 525944 711590
rect 526584 -7654 527224 711590
rect 527864 -7654 528504 711590
rect 529144 -7654 529784 711590
rect 530424 -7654 531064 711590
rect 531704 -7654 532344 711590
rect 532984 -7654 533624 711590
rect 540344 -7654 540984 711590
rect 541624 -7654 542264 711590
rect 542904 -7654 543544 711590
rect 544184 -7654 544824 711590
rect 545464 -7654 546104 711590
rect 546744 -7654 547384 711590
rect 548024 -7654 548664 711590
rect 549304 -7654 549944 711590
rect 556664 -7654 557304 711590
rect 557944 -7654 558584 711590
rect 559224 -7654 559864 711590
rect 560504 -7654 561144 711590
rect 561784 -7654 562424 711590
rect 563064 -7654 563704 711590
rect 564344 -7654 564984 711590
rect 565624 -7654 566264 711590
rect 572984 -7654 573624 711590
rect 574264 -7654 574904 711590
rect 575544 -7654 576184 711590
rect 576824 -7654 577464 711590
rect 578104 -7654 578744 711590
rect 579384 -7654 580024 711590
rect 580664 -7654 581304 711590
rect 581944 -7654 582584 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 6048 151177 6824 161808
rect 7624 151177 8104 161808
rect 8904 151177 9384 161808
rect 10184 151177 10664 161808
rect 11464 151177 18024 161808
rect 18824 151177 19304 161808
rect 20104 151177 20584 161808
rect 21384 151177 23144 161808
rect 23944 151177 24424 161808
rect 25224 151177 25704 161808
rect 26504 151177 26984 161808
rect 27784 151177 34344 161808
rect 35144 151177 35624 161808
rect 36424 151177 36904 161808
rect 37704 151177 39464 161808
rect 40264 151177 40744 161808
rect 41544 151177 42024 161808
rect 42824 151177 43304 161808
rect 44104 151177 50664 161808
rect 51464 151177 51944 161808
rect 52744 151177 53224 161808
rect 54024 151177 55784 161808
rect 56584 151177 57064 161808
rect 57864 151177 58344 161808
rect 59144 151177 59624 161808
rect 60424 151177 66984 161808
rect 67784 151177 68264 161808
rect 69064 151177 69544 161808
rect 70344 151177 72104 161808
rect 72904 151177 73384 161808
rect 74184 151177 74664 161808
rect 75464 151177 75944 161808
rect 76744 151177 83304 161808
rect 84104 151177 84584 161808
rect 85384 151177 85864 161808
rect 86664 151177 88424 161808
rect 89224 151177 89704 161808
rect 90504 151177 90984 161808
rect 91784 151177 92264 161808
rect 93064 151177 99624 161808
rect 100424 151177 100904 161808
rect 101704 151177 102184 161808
rect 102984 151177 104744 161808
rect 105544 151177 106024 161808
rect 106824 151177 107304 161808
rect 108104 151177 108584 161808
rect 109384 151177 115944 161808
rect 116744 151177 117224 161808
rect 118024 151177 118504 161808
rect 119304 151177 121064 161808
rect 121864 151177 122344 161808
rect 123144 151177 123624 161808
rect 124424 151177 124904 161808
rect 125704 151177 132264 161808
rect 133064 151177 133544 161808
rect 134344 151177 134824 161808
rect 135624 151177 137384 161808
rect 138184 151177 138664 161808
rect 139464 151177 139944 161808
rect 140744 151177 141224 161808
rect 142024 151177 148584 161808
rect 149384 151177 149864 161808
rect 150664 151177 151144 161808
rect 151944 151177 153704 161808
rect 154504 151177 154984 161808
rect 155784 151177 156264 161808
rect 157064 151177 157544 161808
rect 158344 151177 162941 161808
rect 6048 4715 162941 151177
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 697256 592650 697896
rect -8726 695976 592650 696616
rect -8726 694696 592650 695336
rect -8726 693416 592650 694056
rect -8726 692136 592650 692776
rect -8726 690856 592650 691496
rect -8726 689576 592650 690216
rect -8726 688296 592650 688936
rect -8726 680936 592650 681576
rect -8726 679656 592650 680296
rect -8726 678376 592650 679016
rect -8726 677096 592650 677736
rect -8726 675816 592650 676456
rect -8726 674536 592650 675176
rect -8726 673256 592650 673896
rect -8726 671976 592650 672616
rect -8726 664616 592650 665256
rect -8726 663336 592650 663976
rect -8726 662056 592650 662696
rect -8726 660776 592650 661416
rect -8726 659496 592650 660136
rect -8726 658216 592650 658856
rect -8726 656936 592650 657576
rect -8726 655656 592650 656296
rect -8726 648296 592650 648936
rect -8726 647016 592650 647656
rect -8726 645736 592650 646376
rect -8726 644456 592650 645096
rect -8726 643176 592650 643816
rect -8726 641896 592650 642536
rect -8726 640616 592650 641256
rect -8726 639336 592650 639976
rect -8726 631976 592650 632616
rect -8726 630696 592650 631336
rect -8726 629416 592650 630056
rect -8726 628136 592650 628776
rect -8726 626856 592650 627496
rect -8726 625576 592650 626216
rect -8726 624296 592650 624936
rect -8726 623016 592650 623656
rect -8726 615656 592650 616296
rect -8726 614376 592650 615016
rect -8726 613096 592650 613736
rect -8726 611816 592650 612456
rect -8726 610536 592650 611176
rect -8726 609256 592650 609896
rect -8726 607976 592650 608616
rect -8726 606696 592650 607336
rect -8726 599336 592650 599976
rect -8726 598056 592650 598696
rect -8726 596776 592650 597416
rect -8726 595496 592650 596136
rect -8726 594216 592650 594856
rect -8726 592936 592650 593576
rect -8726 591656 592650 592296
rect -8726 590376 592650 591016
rect -8726 583016 592650 583656
rect -8726 581736 592650 582376
rect -8726 580456 592650 581096
rect -8726 579176 592650 579816
rect -8726 577896 592650 578536
rect -8726 576616 592650 577256
rect -8726 575336 592650 575976
rect -8726 574056 592650 574696
rect -8726 566696 592650 567336
rect -8726 565416 592650 566056
rect -8726 564136 592650 564776
rect -8726 562856 592650 563496
rect -8726 561576 592650 562216
rect -8726 560296 592650 560936
rect -8726 559016 592650 559656
rect -8726 557736 592650 558376
rect -8726 550376 592650 551016
rect -8726 549096 592650 549736
rect -8726 547816 592650 548456
rect -8726 546536 592650 547176
rect -8726 545256 592650 545896
rect -8726 543976 592650 544616
rect -8726 542696 592650 543336
rect -8726 541416 592650 542056
rect -8726 534056 592650 534696
rect -8726 532776 592650 533416
rect -8726 531496 592650 532136
rect -8726 530216 592650 530856
rect -8726 528936 592650 529576
rect -8726 527656 592650 528296
rect -8726 526376 592650 527016
rect -8726 525096 592650 525736
rect -8726 517736 592650 518376
rect -8726 516456 592650 517096
rect -8726 515176 592650 515816
rect -8726 513896 592650 514536
rect -8726 512616 592650 513256
rect -8726 511336 592650 511976
rect -8726 510056 592650 510696
rect -8726 508776 592650 509416
rect -8726 501416 592650 502056
rect -8726 500136 592650 500776
rect -8726 498856 592650 499496
rect -8726 497576 592650 498216
rect -8726 496296 592650 496936
rect -8726 495016 592650 495656
rect -8726 493736 592650 494376
rect -8726 492456 592650 493096
rect -8726 485096 592650 485736
rect -8726 483816 592650 484456
rect -8726 482536 592650 483176
rect -8726 481256 592650 481896
rect -8726 479976 592650 480616
rect -8726 478696 592650 479336
rect -8726 477416 592650 478056
rect -8726 476136 592650 476776
rect -8726 468776 592650 469416
rect -8726 467496 592650 468136
rect -8726 466216 592650 466856
rect -8726 464936 592650 465576
rect -8726 463656 592650 464296
rect -8726 462376 592650 463016
rect -8726 461096 592650 461736
rect -8726 459816 592650 460456
rect -8726 452456 592650 453096
rect -8726 451176 592650 451816
rect -8726 449896 592650 450536
rect -8726 448616 592650 449256
rect -8726 447336 592650 447976
rect -8726 446056 592650 446696
rect -8726 444776 592650 445416
rect -8726 443496 592650 444136
rect -8726 436136 592650 436776
rect -8726 434856 592650 435496
rect -8726 433576 592650 434216
rect -8726 432296 592650 432936
rect -8726 431016 592650 431656
rect -8726 429736 592650 430376
rect -8726 428456 592650 429096
rect -8726 427176 592650 427816
rect -8726 419816 592650 420456
rect -8726 418536 592650 419176
rect -8726 417256 592650 417896
rect -8726 415976 592650 416616
rect -8726 414696 592650 415336
rect -8726 413416 592650 414056
rect -8726 412136 592650 412776
rect -8726 410856 592650 411496
rect -8726 403496 592650 404136
rect -8726 402216 592650 402856
rect -8726 400936 592650 401576
rect -8726 399656 592650 400296
rect -8726 398376 592650 399016
rect -8726 397096 592650 397736
rect -8726 395816 592650 396456
rect -8726 394536 592650 395176
rect -8726 387176 592650 387816
rect -8726 385896 592650 386536
rect -8726 384616 592650 385256
rect -8726 383336 592650 383976
rect -8726 382056 592650 382696
rect -8726 380776 592650 381416
rect -8726 379496 592650 380136
rect -8726 378216 592650 378856
rect -8726 370856 592650 371496
rect -8726 369576 592650 370216
rect -8726 368296 592650 368936
rect -8726 367016 592650 367656
rect -8726 365736 592650 366376
rect -8726 364456 592650 365096
rect -8726 363176 592650 363816
rect -8726 361896 592650 362536
rect -8726 354536 592650 355176
rect -8726 353256 592650 353896
rect -8726 351976 592650 352616
rect -8726 350696 592650 351336
rect -8726 349416 592650 350056
rect -8726 348136 592650 348776
rect -8726 346856 592650 347496
rect -8726 345576 592650 346216
rect -8726 338216 592650 338856
rect -8726 336936 592650 337576
rect -8726 335656 592650 336296
rect -8726 334376 592650 335016
rect -8726 333096 592650 333736
rect -8726 331816 592650 332456
rect -8726 330536 592650 331176
rect -8726 329256 592650 329896
rect -8726 321896 592650 322536
rect -8726 320616 592650 321256
rect -8726 319336 592650 319976
rect -8726 318056 592650 318696
rect -8726 316776 592650 317416
rect -8726 315496 592650 316136
rect -8726 314216 592650 314856
rect -8726 312936 592650 313576
rect -8726 305576 592650 306216
rect -8726 304296 592650 304936
rect -8726 303016 592650 303656
rect -8726 301736 592650 302376
rect -8726 300456 592650 301096
rect -8726 299176 592650 299816
rect -8726 297896 592650 298536
rect -8726 296616 592650 297256
rect -8726 289256 592650 289896
rect -8726 287976 592650 288616
rect -8726 286696 592650 287336
rect -8726 285416 592650 286056
rect -8726 284136 592650 284776
rect -8726 282856 592650 283496
rect -8726 281576 592650 282216
rect -8726 280296 592650 280936
rect -8726 272936 592650 273576
rect -8726 271656 592650 272296
rect -8726 270376 592650 271016
rect -8726 269096 592650 269736
rect -8726 267816 592650 268456
rect -8726 266536 592650 267176
rect -8726 265256 592650 265896
rect -8726 263976 592650 264616
rect -8726 256616 592650 257256
rect -8726 255336 592650 255976
rect -8726 254056 592650 254696
rect -8726 252776 592650 253416
rect -8726 251496 592650 252136
rect -8726 250216 592650 250856
rect -8726 248936 592650 249576
rect -8726 247656 592650 248296
rect -8726 240296 592650 240936
rect -8726 239016 592650 239656
rect -8726 237736 592650 238376
rect -8726 236456 592650 237096
rect -8726 235176 592650 235816
rect -8726 233896 592650 234536
rect -8726 232616 592650 233256
rect -8726 231336 592650 231976
rect -8726 223976 592650 224616
rect -8726 222696 592650 223336
rect -8726 221416 592650 222056
rect -8726 220136 592650 220776
rect -8726 218856 592650 219496
rect -8726 217576 592650 218216
rect -8726 216296 592650 216936
rect -8726 215016 592650 215656
rect -8726 207656 592650 208296
rect -8726 206376 592650 207016
rect -8726 205096 592650 205736
rect -8726 203816 592650 204456
rect -8726 202536 592650 203176
rect -8726 201256 592650 201896
rect -8726 199976 592650 200616
rect -8726 198696 592650 199336
rect -8726 191336 592650 191976
rect -8726 190056 592650 190696
rect -8726 188776 592650 189416
rect -8726 187496 592650 188136
rect -8726 186216 592650 186856
rect -8726 184936 592650 185576
rect -8726 183656 592650 184296
rect -8726 182376 592650 183016
rect -8726 175016 592650 175656
rect -8726 173736 592650 174376
rect -8726 172456 592650 173096
rect -8726 171176 592650 171816
rect -8726 169896 592650 170536
rect -8726 168616 592650 169256
rect -8726 167336 592650 167976
rect -8726 166056 592650 166696
rect -8726 158696 592650 159336
rect -8726 157416 592650 158056
rect -8726 156136 592650 156776
rect -8726 154856 592650 155496
rect -8726 153576 592650 154216
rect -8726 152296 592650 152936
rect -8726 151016 592650 151656
rect -8726 149736 592650 150376
rect -8726 142376 592650 143016
rect -8726 141096 592650 141736
rect -8726 139816 592650 140456
rect -8726 138536 592650 139176
rect -8726 137256 592650 137896
rect -8726 135976 592650 136616
rect -8726 134696 592650 135336
rect -8726 133416 592650 134056
rect -8726 126056 592650 126696
rect -8726 124776 592650 125416
rect -8726 123496 592650 124136
rect -8726 122216 592650 122856
rect -8726 120936 592650 121576
rect -8726 119656 592650 120296
rect -8726 118376 592650 119016
rect -8726 117096 592650 117736
rect -8726 109736 592650 110376
rect -8726 108456 592650 109096
rect -8726 107176 592650 107816
rect -8726 105896 592650 106536
rect -8726 104616 592650 105256
rect -8726 103336 592650 103976
rect -8726 102056 592650 102696
rect -8726 100776 592650 101416
rect -8726 93416 592650 94056
rect -8726 92136 592650 92776
rect -8726 90856 592650 91496
rect -8726 89576 592650 90216
rect -8726 88296 592650 88936
rect -8726 87016 592650 87656
rect -8726 85736 592650 86376
rect -8726 84456 592650 85096
rect -8726 77096 592650 77736
rect -8726 75816 592650 76456
rect -8726 74536 592650 75176
rect -8726 73256 592650 73896
rect -8726 71976 592650 72616
rect -8726 70696 592650 71336
rect -8726 69416 592650 70056
rect -8726 68136 592650 68776
rect -8726 60776 592650 61416
rect -8726 59496 592650 60136
rect -8726 58216 592650 58856
rect -8726 56936 592650 57576
rect -8726 55656 592650 56296
rect -8726 54376 592650 55016
rect -8726 53096 592650 53736
rect -8726 51816 592650 52456
rect -8726 44456 592650 45096
rect -8726 43176 592650 43816
rect -8726 41896 592650 42536
rect -8726 40616 592650 41256
rect -8726 39336 592650 39976
rect -8726 38056 592650 38696
rect -8726 36776 592650 37416
rect -8726 35496 592650 36136
rect -8726 28136 592650 28776
rect -8726 26856 592650 27496
rect -8726 25576 592650 26216
rect -8726 24296 592650 24936
rect -8726 23016 592650 23656
rect -8726 21736 592650 22376
rect -8726 20456 592650 21096
rect -8726 19176 592650 19816
rect -8726 11816 592650 12456
rect -8726 10536 592650 11176
rect -8726 9256 592650 9896
rect -8726 7976 592650 8616
rect -8726 6696 592650 7336
rect -8726 5416 592650 6056
rect -8726 4136 592650 4776
rect -8726 2856 592650 3496
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew
rlabel metal5 s -8726 688296 592650 688936 6 vccd1
port 532 nsew
rlabel metal5 s -8726 671976 592650 672616 6 vccd1
port 532 nsew
rlabel metal5 s -8726 655656 592650 656296 6 vccd1
port 532 nsew
rlabel metal5 s -8726 639336 592650 639976 6 vccd1
port 532 nsew
rlabel metal5 s -8726 623016 592650 623656 6 vccd1
port 532 nsew
rlabel metal5 s -8726 606696 592650 607336 6 vccd1
port 532 nsew
rlabel metal5 s -8726 590376 592650 591016 6 vccd1
port 532 nsew
rlabel metal5 s -8726 574056 592650 574696 6 vccd1
port 532 nsew
rlabel metal5 s -8726 557736 592650 558376 6 vccd1
port 532 nsew
rlabel metal5 s -8726 541416 592650 542056 6 vccd1
port 532 nsew
rlabel metal5 s -8726 525096 592650 525736 6 vccd1
port 532 nsew
rlabel metal5 s -8726 508776 592650 509416 6 vccd1
port 532 nsew
rlabel metal5 s -8726 492456 592650 493096 6 vccd1
port 532 nsew
rlabel metal5 s -8726 476136 592650 476776 6 vccd1
port 532 nsew
rlabel metal5 s -8726 459816 592650 460456 6 vccd1
port 532 nsew
rlabel metal5 s -8726 443496 592650 444136 6 vccd1
port 532 nsew
rlabel metal5 s -8726 427176 592650 427816 6 vccd1
port 532 nsew
rlabel metal5 s -8726 410856 592650 411496 6 vccd1
port 532 nsew
rlabel metal5 s -8726 394536 592650 395176 6 vccd1
port 532 nsew
rlabel metal5 s -8726 378216 592650 378856 6 vccd1
port 532 nsew
rlabel metal5 s -8726 361896 592650 362536 6 vccd1
port 532 nsew
rlabel metal5 s -8726 345576 592650 346216 6 vccd1
port 532 nsew
rlabel metal5 s -8726 329256 592650 329896 6 vccd1
port 532 nsew
rlabel metal5 s -8726 312936 592650 313576 6 vccd1
port 532 nsew
rlabel metal5 s -8726 296616 592650 297256 6 vccd1
port 532 nsew
rlabel metal5 s -8726 280296 592650 280936 6 vccd1
port 532 nsew
rlabel metal5 s -8726 263976 592650 264616 6 vccd1
port 532 nsew
rlabel metal5 s -8726 247656 592650 248296 6 vccd1
port 532 nsew
rlabel metal5 s -8726 231336 592650 231976 6 vccd1
port 532 nsew
rlabel metal5 s -8726 215016 592650 215656 6 vccd1
port 532 nsew
rlabel metal5 s -8726 198696 592650 199336 6 vccd1
port 532 nsew
rlabel metal5 s -8726 182376 592650 183016 6 vccd1
port 532 nsew
rlabel metal5 s -8726 166056 592650 166696 6 vccd1
port 532 nsew
rlabel metal5 s -8726 149736 592650 150376 6 vccd1
port 532 nsew
rlabel metal5 s -8726 133416 592650 134056 6 vccd1
port 532 nsew
rlabel metal5 s -8726 117096 592650 117736 6 vccd1
port 532 nsew
rlabel metal5 s -8726 100776 592650 101416 6 vccd1
port 532 nsew
rlabel metal5 s -8726 84456 592650 85096 6 vccd1
port 532 nsew
rlabel metal5 s -8726 68136 592650 68776 6 vccd1
port 532 nsew
rlabel metal5 s -8726 51816 592650 52456 6 vccd1
port 532 nsew
rlabel metal5 s -8726 35496 592650 36136 6 vccd1
port 532 nsew
rlabel metal5 s -8726 19176 592650 19816 6 vccd1
port 532 nsew
rlabel metal5 s -8726 2856 592650 3496 6 vccd1
port 532 nsew
rlabel metal4 s 572984 -7654 573624 711590 6 vccd1
port 532 nsew
rlabel metal4 s 556664 -7654 557304 711590 6 vccd1
port 532 nsew
rlabel metal4 s 540344 -7654 540984 711590 6 vccd1
port 532 nsew
rlabel metal4 s 524024 -7654 524664 711590 6 vccd1
port 532 nsew
rlabel metal4 s 507704 -7654 508344 711590 6 vccd1
port 532 nsew
rlabel metal4 s 491384 -7654 492024 711590 6 vccd1
port 532 nsew
rlabel metal4 s 475064 -7654 475704 711590 6 vccd1
port 532 nsew
rlabel metal4 s 458744 -7654 459384 711590 6 vccd1
port 532 nsew
rlabel metal4 s 442424 -7654 443064 711590 6 vccd1
port 532 nsew
rlabel metal4 s 426104 -7654 426744 711590 6 vccd1
port 532 nsew
rlabel metal4 s 409784 -7654 410424 711590 6 vccd1
port 532 nsew
rlabel metal4 s 393464 -7654 394104 711590 6 vccd1
port 532 nsew
rlabel metal4 s 377144 -7654 377784 711590 6 vccd1
port 532 nsew
rlabel metal4 s 360824 -7654 361464 711590 6 vccd1
port 532 nsew
rlabel metal4 s 344504 -7654 345144 711590 6 vccd1
port 532 nsew
rlabel metal4 s 328184 -7654 328824 711590 6 vccd1
port 532 nsew
rlabel metal4 s 311864 -7654 312504 711590 6 vccd1
port 532 nsew
rlabel metal4 s 295544 -7654 296184 711590 6 vccd1
port 532 nsew
rlabel metal4 s 279224 -7654 279864 711590 6 vccd1
port 532 nsew
rlabel metal4 s 262904 -7654 263544 711590 6 vccd1
port 532 nsew
rlabel metal4 s 246584 -7654 247224 711590 6 vccd1
port 532 nsew
rlabel metal4 s 230264 -7654 230904 711590 6 vccd1
port 532 nsew
rlabel metal4 s 213944 -7654 214584 711590 6 vccd1
port 532 nsew
rlabel metal4 s 197624 -7654 198264 711590 6 vccd1
port 532 nsew
rlabel metal4 s 181304 -7654 181944 711590 6 vccd1
port 532 nsew
rlabel metal4 s 164984 151257 165624 711590 6 vccd1
port 532 nsew
rlabel metal4 s 164984 -7654 165624 4575 8 vccd1
port 532 nsew
rlabel metal4 s 148664 151257 149304 711590 6 vccd1
port 532 nsew
rlabel metal4 s 148664 -7654 149304 4575 8 vccd1
port 532 nsew
rlabel metal4 s 132344 151257 132984 711590 6 vccd1
port 532 nsew
rlabel metal4 s 132344 -7654 132984 4575 8 vccd1
port 532 nsew
rlabel metal4 s 116024 151257 116664 711590 6 vccd1
port 532 nsew
rlabel metal4 s 116024 -7654 116664 4575 8 vccd1
port 532 nsew
rlabel metal4 s 99704 151257 100344 711590 6 vccd1
port 532 nsew
rlabel metal4 s 99704 -7654 100344 4575 8 vccd1
port 532 nsew
rlabel metal4 s 83384 151257 84024 711590 6 vccd1
port 532 nsew
rlabel metal4 s 83384 -7654 84024 4575 8 vccd1
port 532 nsew
rlabel metal4 s 67064 151257 67704 711590 6 vccd1
port 532 nsew
rlabel metal4 s 67064 -7654 67704 4575 8 vccd1
port 532 nsew
rlabel metal4 s 50744 151257 51384 711590 6 vccd1
port 532 nsew
rlabel metal4 s 50744 -7654 51384 4575 8 vccd1
port 532 nsew
rlabel metal4 s 34424 151257 35064 711590 6 vccd1
port 532 nsew
rlabel metal4 s 34424 -7654 35064 4575 8 vccd1
port 532 nsew
rlabel metal4 s 18104 151257 18744 711590 6 vccd1
port 532 nsew
rlabel metal4 s 18104 -7654 18744 4575 8 vccd1
port 532 nsew
rlabel metal4 s 1784 -7654 2424 711590 6 vccd1
port 532 nsew
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew
rlabel metal5 s -8726 690856 592650 691496 6 vccd2
port 533 nsew
rlabel metal5 s -8726 674536 592650 675176 6 vccd2
port 533 nsew
rlabel metal5 s -8726 658216 592650 658856 6 vccd2
port 533 nsew
rlabel metal5 s -8726 641896 592650 642536 6 vccd2
port 533 nsew
rlabel metal5 s -8726 625576 592650 626216 6 vccd2
port 533 nsew
rlabel metal5 s -8726 609256 592650 609896 6 vccd2
port 533 nsew
rlabel metal5 s -8726 592936 592650 593576 6 vccd2
port 533 nsew
rlabel metal5 s -8726 576616 592650 577256 6 vccd2
port 533 nsew
rlabel metal5 s -8726 560296 592650 560936 6 vccd2
port 533 nsew
rlabel metal5 s -8726 543976 592650 544616 6 vccd2
port 533 nsew
rlabel metal5 s -8726 527656 592650 528296 6 vccd2
port 533 nsew
rlabel metal5 s -8726 511336 592650 511976 6 vccd2
port 533 nsew
rlabel metal5 s -8726 495016 592650 495656 6 vccd2
port 533 nsew
rlabel metal5 s -8726 478696 592650 479336 6 vccd2
port 533 nsew
rlabel metal5 s -8726 462376 592650 463016 6 vccd2
port 533 nsew
rlabel metal5 s -8726 446056 592650 446696 6 vccd2
port 533 nsew
rlabel metal5 s -8726 429736 592650 430376 6 vccd2
port 533 nsew
rlabel metal5 s -8726 413416 592650 414056 6 vccd2
port 533 nsew
rlabel metal5 s -8726 397096 592650 397736 6 vccd2
port 533 nsew
rlabel metal5 s -8726 380776 592650 381416 6 vccd2
port 533 nsew
rlabel metal5 s -8726 364456 592650 365096 6 vccd2
port 533 nsew
rlabel metal5 s -8726 348136 592650 348776 6 vccd2
port 533 nsew
rlabel metal5 s -8726 331816 592650 332456 6 vccd2
port 533 nsew
rlabel metal5 s -8726 315496 592650 316136 6 vccd2
port 533 nsew
rlabel metal5 s -8726 299176 592650 299816 6 vccd2
port 533 nsew
rlabel metal5 s -8726 282856 592650 283496 6 vccd2
port 533 nsew
rlabel metal5 s -8726 266536 592650 267176 6 vccd2
port 533 nsew
rlabel metal5 s -8726 250216 592650 250856 6 vccd2
port 533 nsew
rlabel metal5 s -8726 233896 592650 234536 6 vccd2
port 533 nsew
rlabel metal5 s -8726 217576 592650 218216 6 vccd2
port 533 nsew
rlabel metal5 s -8726 201256 592650 201896 6 vccd2
port 533 nsew
rlabel metal5 s -8726 184936 592650 185576 6 vccd2
port 533 nsew
rlabel metal5 s -8726 168616 592650 169256 6 vccd2
port 533 nsew
rlabel metal5 s -8726 152296 592650 152936 6 vccd2
port 533 nsew
rlabel metal5 s -8726 135976 592650 136616 6 vccd2
port 533 nsew
rlabel metal5 s -8726 119656 592650 120296 6 vccd2
port 533 nsew
rlabel metal5 s -8726 103336 592650 103976 6 vccd2
port 533 nsew
rlabel metal5 s -8726 87016 592650 87656 6 vccd2
port 533 nsew
rlabel metal5 s -8726 70696 592650 71336 6 vccd2
port 533 nsew
rlabel metal5 s -8726 54376 592650 55016 6 vccd2
port 533 nsew
rlabel metal5 s -8726 38056 592650 38696 6 vccd2
port 533 nsew
rlabel metal5 s -8726 21736 592650 22376 6 vccd2
port 533 nsew
rlabel metal5 s -8726 5416 592650 6056 6 vccd2
port 533 nsew
rlabel metal4 s 575544 -7654 576184 711590 6 vccd2
port 533 nsew
rlabel metal4 s 559224 -7654 559864 711590 6 vccd2
port 533 nsew
rlabel metal4 s 542904 -7654 543544 711590 6 vccd2
port 533 nsew
rlabel metal4 s 526584 -7654 527224 711590 6 vccd2
port 533 nsew
rlabel metal4 s 510264 -7654 510904 711590 6 vccd2
port 533 nsew
rlabel metal4 s 493944 -7654 494584 711590 6 vccd2
port 533 nsew
rlabel metal4 s 477624 -7654 478264 711590 6 vccd2
port 533 nsew
rlabel metal4 s 461304 -7654 461944 711590 6 vccd2
port 533 nsew
rlabel metal4 s 444984 -7654 445624 711590 6 vccd2
port 533 nsew
rlabel metal4 s 428664 -7654 429304 711590 6 vccd2
port 533 nsew
rlabel metal4 s 412344 -7654 412984 711590 6 vccd2
port 533 nsew
rlabel metal4 s 396024 -7654 396664 711590 6 vccd2
port 533 nsew
rlabel metal4 s 379704 -7654 380344 711590 6 vccd2
port 533 nsew
rlabel metal4 s 363384 -7654 364024 711590 6 vccd2
port 533 nsew
rlabel metal4 s 347064 -7654 347704 711590 6 vccd2
port 533 nsew
rlabel metal4 s 330744 -7654 331384 711590 6 vccd2
port 533 nsew
rlabel metal4 s 314424 -7654 315064 711590 6 vccd2
port 533 nsew
rlabel metal4 s 298104 -7654 298744 711590 6 vccd2
port 533 nsew
rlabel metal4 s 281784 -7654 282424 711590 6 vccd2
port 533 nsew
rlabel metal4 s 265464 -7654 266104 711590 6 vccd2
port 533 nsew
rlabel metal4 s 249144 -7654 249784 711590 6 vccd2
port 533 nsew
rlabel metal4 s 232824 -7654 233464 711590 6 vccd2
port 533 nsew
rlabel metal4 s 216504 -7654 217144 711590 6 vccd2
port 533 nsew
rlabel metal4 s 200184 -7654 200824 711590 6 vccd2
port 533 nsew
rlabel metal4 s 183864 -7654 184504 711590 6 vccd2
port 533 nsew
rlabel metal4 s 167544 -7654 168184 711590 6 vccd2
port 533 nsew
rlabel metal4 s 151224 151257 151864 711590 6 vccd2
port 533 nsew
rlabel metal4 s 134904 151257 135544 711590 6 vccd2
port 533 nsew
rlabel metal4 s 118584 151257 119224 711590 6 vccd2
port 533 nsew
rlabel metal4 s 102264 151257 102904 711590 6 vccd2
port 533 nsew
rlabel metal4 s 85944 151257 86584 711590 6 vccd2
port 533 nsew
rlabel metal4 s 69624 151257 70264 711590 6 vccd2
port 533 nsew
rlabel metal4 s 53304 151257 53944 711590 6 vccd2
port 533 nsew
rlabel metal4 s 36984 151257 37624 711590 6 vccd2
port 533 nsew
rlabel metal4 s 20664 151257 21304 711590 6 vccd2
port 533 nsew
rlabel metal4 s 4344 -7654 4984 711590 6 vccd2
port 533 nsew
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew
rlabel metal5 s -8726 693416 592650 694056 6 vdda1
port 534 nsew
rlabel metal5 s -8726 677096 592650 677736 6 vdda1
port 534 nsew
rlabel metal5 s -8726 660776 592650 661416 6 vdda1
port 534 nsew
rlabel metal5 s -8726 644456 592650 645096 6 vdda1
port 534 nsew
rlabel metal5 s -8726 628136 592650 628776 6 vdda1
port 534 nsew
rlabel metal5 s -8726 611816 592650 612456 6 vdda1
port 534 nsew
rlabel metal5 s -8726 595496 592650 596136 6 vdda1
port 534 nsew
rlabel metal5 s -8726 579176 592650 579816 6 vdda1
port 534 nsew
rlabel metal5 s -8726 562856 592650 563496 6 vdda1
port 534 nsew
rlabel metal5 s -8726 546536 592650 547176 6 vdda1
port 534 nsew
rlabel metal5 s -8726 530216 592650 530856 6 vdda1
port 534 nsew
rlabel metal5 s -8726 513896 592650 514536 6 vdda1
port 534 nsew
rlabel metal5 s -8726 497576 592650 498216 6 vdda1
port 534 nsew
rlabel metal5 s -8726 481256 592650 481896 6 vdda1
port 534 nsew
rlabel metal5 s -8726 464936 592650 465576 6 vdda1
port 534 nsew
rlabel metal5 s -8726 448616 592650 449256 6 vdda1
port 534 nsew
rlabel metal5 s -8726 432296 592650 432936 6 vdda1
port 534 nsew
rlabel metal5 s -8726 415976 592650 416616 6 vdda1
port 534 nsew
rlabel metal5 s -8726 399656 592650 400296 6 vdda1
port 534 nsew
rlabel metal5 s -8726 383336 592650 383976 6 vdda1
port 534 nsew
rlabel metal5 s -8726 367016 592650 367656 6 vdda1
port 534 nsew
rlabel metal5 s -8726 350696 592650 351336 6 vdda1
port 534 nsew
rlabel metal5 s -8726 334376 592650 335016 6 vdda1
port 534 nsew
rlabel metal5 s -8726 318056 592650 318696 6 vdda1
port 534 nsew
rlabel metal5 s -8726 301736 592650 302376 6 vdda1
port 534 nsew
rlabel metal5 s -8726 285416 592650 286056 6 vdda1
port 534 nsew
rlabel metal5 s -8726 269096 592650 269736 6 vdda1
port 534 nsew
rlabel metal5 s -8726 252776 592650 253416 6 vdda1
port 534 nsew
rlabel metal5 s -8726 236456 592650 237096 6 vdda1
port 534 nsew
rlabel metal5 s -8726 220136 592650 220776 6 vdda1
port 534 nsew
rlabel metal5 s -8726 203816 592650 204456 6 vdda1
port 534 nsew
rlabel metal5 s -8726 187496 592650 188136 6 vdda1
port 534 nsew
rlabel metal5 s -8726 171176 592650 171816 6 vdda1
port 534 nsew
rlabel metal5 s -8726 154856 592650 155496 6 vdda1
port 534 nsew
rlabel metal5 s -8726 138536 592650 139176 6 vdda1
port 534 nsew
rlabel metal5 s -8726 122216 592650 122856 6 vdda1
port 534 nsew
rlabel metal5 s -8726 105896 592650 106536 6 vdda1
port 534 nsew
rlabel metal5 s -8726 89576 592650 90216 6 vdda1
port 534 nsew
rlabel metal5 s -8726 73256 592650 73896 6 vdda1
port 534 nsew
rlabel metal5 s -8726 56936 592650 57576 6 vdda1
port 534 nsew
rlabel metal5 s -8726 40616 592650 41256 6 vdda1
port 534 nsew
rlabel metal5 s -8726 24296 592650 24936 6 vdda1
port 534 nsew
rlabel metal5 s -8726 7976 592650 8616 6 vdda1
port 534 nsew
rlabel metal4 s 578104 -7654 578744 711590 6 vdda1
port 534 nsew
rlabel metal4 s 561784 -7654 562424 711590 6 vdda1
port 534 nsew
rlabel metal4 s 545464 -7654 546104 711590 6 vdda1
port 534 nsew
rlabel metal4 s 529144 -7654 529784 711590 6 vdda1
port 534 nsew
rlabel metal4 s 512824 -7654 513464 711590 6 vdda1
port 534 nsew
rlabel metal4 s 496504 -7654 497144 711590 6 vdda1
port 534 nsew
rlabel metal4 s 480184 -7654 480824 711590 6 vdda1
port 534 nsew
rlabel metal4 s 463864 -7654 464504 711590 6 vdda1
port 534 nsew
rlabel metal4 s 447544 -7654 448184 711590 6 vdda1
port 534 nsew
rlabel metal4 s 431224 -7654 431864 711590 6 vdda1
port 534 nsew
rlabel metal4 s 414904 -7654 415544 711590 6 vdda1
port 534 nsew
rlabel metal4 s 398584 -7654 399224 711590 6 vdda1
port 534 nsew
rlabel metal4 s 382264 -7654 382904 711590 6 vdda1
port 534 nsew
rlabel metal4 s 365944 -7654 366584 711590 6 vdda1
port 534 nsew
rlabel metal4 s 349624 -7654 350264 711590 6 vdda1
port 534 nsew
rlabel metal4 s 333304 -7654 333944 711590 6 vdda1
port 534 nsew
rlabel metal4 s 316984 -7654 317624 711590 6 vdda1
port 534 nsew
rlabel metal4 s 300664 -7654 301304 711590 6 vdda1
port 534 nsew
rlabel metal4 s 284344 -7654 284984 711590 6 vdda1
port 534 nsew
rlabel metal4 s 268024 -7654 268664 711590 6 vdda1
port 534 nsew
rlabel metal4 s 251704 -7654 252344 711590 6 vdda1
port 534 nsew
rlabel metal4 s 235384 -7654 236024 711590 6 vdda1
port 534 nsew
rlabel metal4 s 219064 -7654 219704 711590 6 vdda1
port 534 nsew
rlabel metal4 s 202744 -7654 203384 711590 6 vdda1
port 534 nsew
rlabel metal4 s 186424 -7654 187064 711590 6 vdda1
port 534 nsew
rlabel metal4 s 170104 -7654 170744 711590 6 vdda1
port 534 nsew
rlabel metal4 s 153784 151257 154424 711590 6 vdda1
port 534 nsew
rlabel metal4 s 137464 151257 138104 711590 6 vdda1
port 534 nsew
rlabel metal4 s 121144 151257 121784 711590 6 vdda1
port 534 nsew
rlabel metal4 s 104824 151257 105464 711590 6 vdda1
port 534 nsew
rlabel metal4 s 88504 151257 89144 711590 6 vdda1
port 534 nsew
rlabel metal4 s 72184 151257 72824 711590 6 vdda1
port 534 nsew
rlabel metal4 s 55864 151257 56504 711590 6 vdda1
port 534 nsew
rlabel metal4 s 39544 151257 40184 711590 6 vdda1
port 534 nsew
rlabel metal4 s 23224 151257 23864 711590 6 vdda1
port 534 nsew
rlabel metal4 s 6904 151257 7544 711590 6 vdda1
port 534 nsew
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew
rlabel metal5 s -8726 695976 592650 696616 6 vdda2
port 535 nsew
rlabel metal5 s -8726 679656 592650 680296 6 vdda2
port 535 nsew
rlabel metal5 s -8726 663336 592650 663976 6 vdda2
port 535 nsew
rlabel metal5 s -8726 647016 592650 647656 6 vdda2
port 535 nsew
rlabel metal5 s -8726 630696 592650 631336 6 vdda2
port 535 nsew
rlabel metal5 s -8726 614376 592650 615016 6 vdda2
port 535 nsew
rlabel metal5 s -8726 598056 592650 598696 6 vdda2
port 535 nsew
rlabel metal5 s -8726 581736 592650 582376 6 vdda2
port 535 nsew
rlabel metal5 s -8726 565416 592650 566056 6 vdda2
port 535 nsew
rlabel metal5 s -8726 549096 592650 549736 6 vdda2
port 535 nsew
rlabel metal5 s -8726 532776 592650 533416 6 vdda2
port 535 nsew
rlabel metal5 s -8726 516456 592650 517096 6 vdda2
port 535 nsew
rlabel metal5 s -8726 500136 592650 500776 6 vdda2
port 535 nsew
rlabel metal5 s -8726 483816 592650 484456 6 vdda2
port 535 nsew
rlabel metal5 s -8726 467496 592650 468136 6 vdda2
port 535 nsew
rlabel metal5 s -8726 451176 592650 451816 6 vdda2
port 535 nsew
rlabel metal5 s -8726 434856 592650 435496 6 vdda2
port 535 nsew
rlabel metal5 s -8726 418536 592650 419176 6 vdda2
port 535 nsew
rlabel metal5 s -8726 402216 592650 402856 6 vdda2
port 535 nsew
rlabel metal5 s -8726 385896 592650 386536 6 vdda2
port 535 nsew
rlabel metal5 s -8726 369576 592650 370216 6 vdda2
port 535 nsew
rlabel metal5 s -8726 353256 592650 353896 6 vdda2
port 535 nsew
rlabel metal5 s -8726 336936 592650 337576 6 vdda2
port 535 nsew
rlabel metal5 s -8726 320616 592650 321256 6 vdda2
port 535 nsew
rlabel metal5 s -8726 304296 592650 304936 6 vdda2
port 535 nsew
rlabel metal5 s -8726 287976 592650 288616 6 vdda2
port 535 nsew
rlabel metal5 s -8726 271656 592650 272296 6 vdda2
port 535 nsew
rlabel metal5 s -8726 255336 592650 255976 6 vdda2
port 535 nsew
rlabel metal5 s -8726 239016 592650 239656 6 vdda2
port 535 nsew
rlabel metal5 s -8726 222696 592650 223336 6 vdda2
port 535 nsew
rlabel metal5 s -8726 206376 592650 207016 6 vdda2
port 535 nsew
rlabel metal5 s -8726 190056 592650 190696 6 vdda2
port 535 nsew
rlabel metal5 s -8726 173736 592650 174376 6 vdda2
port 535 nsew
rlabel metal5 s -8726 157416 592650 158056 6 vdda2
port 535 nsew
rlabel metal5 s -8726 141096 592650 141736 6 vdda2
port 535 nsew
rlabel metal5 s -8726 124776 592650 125416 6 vdda2
port 535 nsew
rlabel metal5 s -8726 108456 592650 109096 6 vdda2
port 535 nsew
rlabel metal5 s -8726 92136 592650 92776 6 vdda2
port 535 nsew
rlabel metal5 s -8726 75816 592650 76456 6 vdda2
port 535 nsew
rlabel metal5 s -8726 59496 592650 60136 6 vdda2
port 535 nsew
rlabel metal5 s -8726 43176 592650 43816 6 vdda2
port 535 nsew
rlabel metal5 s -8726 26856 592650 27496 6 vdda2
port 535 nsew
rlabel metal5 s -8726 10536 592650 11176 6 vdda2
port 535 nsew
rlabel metal4 s 580664 -7654 581304 711590 6 vdda2
port 535 nsew
rlabel metal4 s 564344 -7654 564984 711590 6 vdda2
port 535 nsew
rlabel metal4 s 548024 -7654 548664 711590 6 vdda2
port 535 nsew
rlabel metal4 s 531704 -7654 532344 711590 6 vdda2
port 535 nsew
rlabel metal4 s 515384 -7654 516024 711590 6 vdda2
port 535 nsew
rlabel metal4 s 499064 -7654 499704 711590 6 vdda2
port 535 nsew
rlabel metal4 s 482744 -7654 483384 711590 6 vdda2
port 535 nsew
rlabel metal4 s 466424 -7654 467064 711590 6 vdda2
port 535 nsew
rlabel metal4 s 450104 -7654 450744 711590 6 vdda2
port 535 nsew
rlabel metal4 s 433784 -7654 434424 711590 6 vdda2
port 535 nsew
rlabel metal4 s 417464 -7654 418104 711590 6 vdda2
port 535 nsew
rlabel metal4 s 401144 -7654 401784 711590 6 vdda2
port 535 nsew
rlabel metal4 s 384824 -7654 385464 711590 6 vdda2
port 535 nsew
rlabel metal4 s 368504 -7654 369144 711590 6 vdda2
port 535 nsew
rlabel metal4 s 352184 -7654 352824 711590 6 vdda2
port 535 nsew
rlabel metal4 s 335864 -7654 336504 711590 6 vdda2
port 535 nsew
rlabel metal4 s 319544 -7654 320184 711590 6 vdda2
port 535 nsew
rlabel metal4 s 303224 -7654 303864 711590 6 vdda2
port 535 nsew
rlabel metal4 s 286904 -7654 287544 711590 6 vdda2
port 535 nsew
rlabel metal4 s 270584 -7654 271224 711590 6 vdda2
port 535 nsew
rlabel metal4 s 254264 -7654 254904 711590 6 vdda2
port 535 nsew
rlabel metal4 s 237944 -7654 238584 711590 6 vdda2
port 535 nsew
rlabel metal4 s 221624 -7654 222264 711590 6 vdda2
port 535 nsew
rlabel metal4 s 205304 -7654 205944 711590 6 vdda2
port 535 nsew
rlabel metal4 s 188984 -7654 189624 711590 6 vdda2
port 535 nsew
rlabel metal4 s 172664 -7654 173304 711590 6 vdda2
port 535 nsew
rlabel metal4 s 156344 151257 156984 711590 6 vdda2
port 535 nsew
rlabel metal4 s 140024 151257 140664 711590 6 vdda2
port 535 nsew
rlabel metal4 s 123704 151257 124344 711590 6 vdda2
port 535 nsew
rlabel metal4 s 107384 151257 108024 711590 6 vdda2
port 535 nsew
rlabel metal4 s 91064 151257 91704 711590 6 vdda2
port 535 nsew
rlabel metal4 s 74744 151257 75384 711590 6 vdda2
port 535 nsew
rlabel metal4 s 58424 151257 59064 711590 6 vdda2
port 535 nsew
rlabel metal4 s 42104 151257 42744 711590 6 vdda2
port 535 nsew
rlabel metal4 s 25784 151257 26424 711590 6 vdda2
port 535 nsew
rlabel metal4 s 9464 151257 10104 711590 6 vdda2
port 535 nsew
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew
rlabel metal5 s -8726 694696 592650 695336 6 vssa1
port 536 nsew
rlabel metal5 s -8726 678376 592650 679016 6 vssa1
port 536 nsew
rlabel metal5 s -8726 662056 592650 662696 6 vssa1
port 536 nsew
rlabel metal5 s -8726 645736 592650 646376 6 vssa1
port 536 nsew
rlabel metal5 s -8726 629416 592650 630056 6 vssa1
port 536 nsew
rlabel metal5 s -8726 613096 592650 613736 6 vssa1
port 536 nsew
rlabel metal5 s -8726 596776 592650 597416 6 vssa1
port 536 nsew
rlabel metal5 s -8726 580456 592650 581096 6 vssa1
port 536 nsew
rlabel metal5 s -8726 564136 592650 564776 6 vssa1
port 536 nsew
rlabel metal5 s -8726 547816 592650 548456 6 vssa1
port 536 nsew
rlabel metal5 s -8726 531496 592650 532136 6 vssa1
port 536 nsew
rlabel metal5 s -8726 515176 592650 515816 6 vssa1
port 536 nsew
rlabel metal5 s -8726 498856 592650 499496 6 vssa1
port 536 nsew
rlabel metal5 s -8726 482536 592650 483176 6 vssa1
port 536 nsew
rlabel metal5 s -8726 466216 592650 466856 6 vssa1
port 536 nsew
rlabel metal5 s -8726 449896 592650 450536 6 vssa1
port 536 nsew
rlabel metal5 s -8726 433576 592650 434216 6 vssa1
port 536 nsew
rlabel metal5 s -8726 417256 592650 417896 6 vssa1
port 536 nsew
rlabel metal5 s -8726 400936 592650 401576 6 vssa1
port 536 nsew
rlabel metal5 s -8726 384616 592650 385256 6 vssa1
port 536 nsew
rlabel metal5 s -8726 368296 592650 368936 6 vssa1
port 536 nsew
rlabel metal5 s -8726 351976 592650 352616 6 vssa1
port 536 nsew
rlabel metal5 s -8726 335656 592650 336296 6 vssa1
port 536 nsew
rlabel metal5 s -8726 319336 592650 319976 6 vssa1
port 536 nsew
rlabel metal5 s -8726 303016 592650 303656 6 vssa1
port 536 nsew
rlabel metal5 s -8726 286696 592650 287336 6 vssa1
port 536 nsew
rlabel metal5 s -8726 270376 592650 271016 6 vssa1
port 536 nsew
rlabel metal5 s -8726 254056 592650 254696 6 vssa1
port 536 nsew
rlabel metal5 s -8726 237736 592650 238376 6 vssa1
port 536 nsew
rlabel metal5 s -8726 221416 592650 222056 6 vssa1
port 536 nsew
rlabel metal5 s -8726 205096 592650 205736 6 vssa1
port 536 nsew
rlabel metal5 s -8726 188776 592650 189416 6 vssa1
port 536 nsew
rlabel metal5 s -8726 172456 592650 173096 6 vssa1
port 536 nsew
rlabel metal5 s -8726 156136 592650 156776 6 vssa1
port 536 nsew
rlabel metal5 s -8726 139816 592650 140456 6 vssa1
port 536 nsew
rlabel metal5 s -8726 123496 592650 124136 6 vssa1
port 536 nsew
rlabel metal5 s -8726 107176 592650 107816 6 vssa1
port 536 nsew
rlabel metal5 s -8726 90856 592650 91496 6 vssa1
port 536 nsew
rlabel metal5 s -8726 74536 592650 75176 6 vssa1
port 536 nsew
rlabel metal5 s -8726 58216 592650 58856 6 vssa1
port 536 nsew
rlabel metal5 s -8726 41896 592650 42536 6 vssa1
port 536 nsew
rlabel metal5 s -8726 25576 592650 26216 6 vssa1
port 536 nsew
rlabel metal5 s -8726 9256 592650 9896 6 vssa1
port 536 nsew
rlabel metal4 s 579384 -7654 580024 711590 6 vssa1
port 536 nsew
rlabel metal4 s 563064 -7654 563704 711590 6 vssa1
port 536 nsew
rlabel metal4 s 546744 -7654 547384 711590 6 vssa1
port 536 nsew
rlabel metal4 s 530424 -7654 531064 711590 6 vssa1
port 536 nsew
rlabel metal4 s 514104 -7654 514744 711590 6 vssa1
port 536 nsew
rlabel metal4 s 497784 -7654 498424 711590 6 vssa1
port 536 nsew
rlabel metal4 s 481464 -7654 482104 711590 6 vssa1
port 536 nsew
rlabel metal4 s 465144 -7654 465784 711590 6 vssa1
port 536 nsew
rlabel metal4 s 448824 -7654 449464 711590 6 vssa1
port 536 nsew
rlabel metal4 s 432504 -7654 433144 711590 6 vssa1
port 536 nsew
rlabel metal4 s 416184 -7654 416824 711590 6 vssa1
port 536 nsew
rlabel metal4 s 399864 -7654 400504 711590 6 vssa1
port 536 nsew
rlabel metal4 s 383544 -7654 384184 711590 6 vssa1
port 536 nsew
rlabel metal4 s 367224 -7654 367864 711590 6 vssa1
port 536 nsew
rlabel metal4 s 350904 -7654 351544 711590 6 vssa1
port 536 nsew
rlabel metal4 s 334584 -7654 335224 711590 6 vssa1
port 536 nsew
rlabel metal4 s 318264 -7654 318904 711590 6 vssa1
port 536 nsew
rlabel metal4 s 301944 -7654 302584 711590 6 vssa1
port 536 nsew
rlabel metal4 s 285624 -7654 286264 711590 6 vssa1
port 536 nsew
rlabel metal4 s 269304 -7654 269944 711590 6 vssa1
port 536 nsew
rlabel metal4 s 252984 -7654 253624 711590 6 vssa1
port 536 nsew
rlabel metal4 s 236664 -7654 237304 711590 6 vssa1
port 536 nsew
rlabel metal4 s 220344 -7654 220984 711590 6 vssa1
port 536 nsew
rlabel metal4 s 204024 -7654 204664 711590 6 vssa1
port 536 nsew
rlabel metal4 s 187704 -7654 188344 711590 6 vssa1
port 536 nsew
rlabel metal4 s 171384 -7654 172024 711590 6 vssa1
port 536 nsew
rlabel metal4 s 155064 151257 155704 711590 6 vssa1
port 536 nsew
rlabel metal4 s 138744 151257 139384 711590 6 vssa1
port 536 nsew
rlabel metal4 s 122424 151257 123064 711590 6 vssa1
port 536 nsew
rlabel metal4 s 106104 151257 106744 711590 6 vssa1
port 536 nsew
rlabel metal4 s 89784 151257 90424 711590 6 vssa1
port 536 nsew
rlabel metal4 s 73464 151257 74104 711590 6 vssa1
port 536 nsew
rlabel metal4 s 57144 151257 57784 711590 6 vssa1
port 536 nsew
rlabel metal4 s 40824 151257 41464 711590 6 vssa1
port 536 nsew
rlabel metal4 s 24504 151257 25144 711590 6 vssa1
port 536 nsew
rlabel metal4 s 8184 151257 8824 711590 6 vssa1
port 536 nsew
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew
rlabel metal5 s -8726 697256 592650 697896 6 vssa2
port 537 nsew
rlabel metal5 s -8726 680936 592650 681576 6 vssa2
port 537 nsew
rlabel metal5 s -8726 664616 592650 665256 6 vssa2
port 537 nsew
rlabel metal5 s -8726 648296 592650 648936 6 vssa2
port 537 nsew
rlabel metal5 s -8726 631976 592650 632616 6 vssa2
port 537 nsew
rlabel metal5 s -8726 615656 592650 616296 6 vssa2
port 537 nsew
rlabel metal5 s -8726 599336 592650 599976 6 vssa2
port 537 nsew
rlabel metal5 s -8726 583016 592650 583656 6 vssa2
port 537 nsew
rlabel metal5 s -8726 566696 592650 567336 6 vssa2
port 537 nsew
rlabel metal5 s -8726 550376 592650 551016 6 vssa2
port 537 nsew
rlabel metal5 s -8726 534056 592650 534696 6 vssa2
port 537 nsew
rlabel metal5 s -8726 517736 592650 518376 6 vssa2
port 537 nsew
rlabel metal5 s -8726 501416 592650 502056 6 vssa2
port 537 nsew
rlabel metal5 s -8726 485096 592650 485736 6 vssa2
port 537 nsew
rlabel metal5 s -8726 468776 592650 469416 6 vssa2
port 537 nsew
rlabel metal5 s -8726 452456 592650 453096 6 vssa2
port 537 nsew
rlabel metal5 s -8726 436136 592650 436776 6 vssa2
port 537 nsew
rlabel metal5 s -8726 419816 592650 420456 6 vssa2
port 537 nsew
rlabel metal5 s -8726 403496 592650 404136 6 vssa2
port 537 nsew
rlabel metal5 s -8726 387176 592650 387816 6 vssa2
port 537 nsew
rlabel metal5 s -8726 370856 592650 371496 6 vssa2
port 537 nsew
rlabel metal5 s -8726 354536 592650 355176 6 vssa2
port 537 nsew
rlabel metal5 s -8726 338216 592650 338856 6 vssa2
port 537 nsew
rlabel metal5 s -8726 321896 592650 322536 6 vssa2
port 537 nsew
rlabel metal5 s -8726 305576 592650 306216 6 vssa2
port 537 nsew
rlabel metal5 s -8726 289256 592650 289896 6 vssa2
port 537 nsew
rlabel metal5 s -8726 272936 592650 273576 6 vssa2
port 537 nsew
rlabel metal5 s -8726 256616 592650 257256 6 vssa2
port 537 nsew
rlabel metal5 s -8726 240296 592650 240936 6 vssa2
port 537 nsew
rlabel metal5 s -8726 223976 592650 224616 6 vssa2
port 537 nsew
rlabel metal5 s -8726 207656 592650 208296 6 vssa2
port 537 nsew
rlabel metal5 s -8726 191336 592650 191976 6 vssa2
port 537 nsew
rlabel metal5 s -8726 175016 592650 175656 6 vssa2
port 537 nsew
rlabel metal5 s -8726 158696 592650 159336 6 vssa2
port 537 nsew
rlabel metal5 s -8726 142376 592650 143016 6 vssa2
port 537 nsew
rlabel metal5 s -8726 126056 592650 126696 6 vssa2
port 537 nsew
rlabel metal5 s -8726 109736 592650 110376 6 vssa2
port 537 nsew
rlabel metal5 s -8726 93416 592650 94056 6 vssa2
port 537 nsew
rlabel metal5 s -8726 77096 592650 77736 6 vssa2
port 537 nsew
rlabel metal5 s -8726 60776 592650 61416 6 vssa2
port 537 nsew
rlabel metal5 s -8726 44456 592650 45096 6 vssa2
port 537 nsew
rlabel metal5 s -8726 28136 592650 28776 6 vssa2
port 537 nsew
rlabel metal5 s -8726 11816 592650 12456 6 vssa2
port 537 nsew
rlabel metal4 s 581944 -7654 582584 711590 6 vssa2
port 537 nsew
rlabel metal4 s 565624 -7654 566264 711590 6 vssa2
port 537 nsew
rlabel metal4 s 549304 -7654 549944 711590 6 vssa2
port 537 nsew
rlabel metal4 s 532984 -7654 533624 711590 6 vssa2
port 537 nsew
rlabel metal4 s 516664 -7654 517304 711590 6 vssa2
port 537 nsew
rlabel metal4 s 500344 -7654 500984 711590 6 vssa2
port 537 nsew
rlabel metal4 s 484024 -7654 484664 711590 6 vssa2
port 537 nsew
rlabel metal4 s 467704 -7654 468344 711590 6 vssa2
port 537 nsew
rlabel metal4 s 451384 -7654 452024 711590 6 vssa2
port 537 nsew
rlabel metal4 s 435064 -7654 435704 711590 6 vssa2
port 537 nsew
rlabel metal4 s 418744 -7654 419384 711590 6 vssa2
port 537 nsew
rlabel metal4 s 402424 -7654 403064 711590 6 vssa2
port 537 nsew
rlabel metal4 s 386104 -7654 386744 711590 6 vssa2
port 537 nsew
rlabel metal4 s 369784 -7654 370424 711590 6 vssa2
port 537 nsew
rlabel metal4 s 353464 -7654 354104 711590 6 vssa2
port 537 nsew
rlabel metal4 s 337144 -7654 337784 711590 6 vssa2
port 537 nsew
rlabel metal4 s 320824 -7654 321464 711590 6 vssa2
port 537 nsew
rlabel metal4 s 304504 -7654 305144 711590 6 vssa2
port 537 nsew
rlabel metal4 s 288184 -7654 288824 711590 6 vssa2
port 537 nsew
rlabel metal4 s 271864 -7654 272504 711590 6 vssa2
port 537 nsew
rlabel metal4 s 255544 -7654 256184 711590 6 vssa2
port 537 nsew
rlabel metal4 s 239224 -7654 239864 711590 6 vssa2
port 537 nsew
rlabel metal4 s 222904 -7654 223544 711590 6 vssa2
port 537 nsew
rlabel metal4 s 206584 -7654 207224 711590 6 vssa2
port 537 nsew
rlabel metal4 s 190264 -7654 190904 711590 6 vssa2
port 537 nsew
rlabel metal4 s 173944 -7654 174584 711590 6 vssa2
port 537 nsew
rlabel metal4 s 157624 151257 158264 711590 6 vssa2
port 537 nsew
rlabel metal4 s 141304 151257 141944 711590 6 vssa2
port 537 nsew
rlabel metal4 s 124984 151257 125624 711590 6 vssa2
port 537 nsew
rlabel metal4 s 108664 151257 109304 711590 6 vssa2
port 537 nsew
rlabel metal4 s 92344 151257 92984 711590 6 vssa2
port 537 nsew
rlabel metal4 s 76024 151257 76664 711590 6 vssa2
port 537 nsew
rlabel metal4 s 59704 151257 60344 711590 6 vssa2
port 537 nsew
rlabel metal4 s 43384 151257 44024 711590 6 vssa2
port 537 nsew
rlabel metal4 s 27064 151257 27704 711590 6 vssa2
port 537 nsew
rlabel metal4 s 10744 151257 11384 711590 6 vssa2
port 537 nsew
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew
rlabel metal5 s -8726 689576 592650 690216 6 vssd1
port 538 nsew
rlabel metal5 s -8726 673256 592650 673896 6 vssd1
port 538 nsew
rlabel metal5 s -8726 656936 592650 657576 6 vssd1
port 538 nsew
rlabel metal5 s -8726 640616 592650 641256 6 vssd1
port 538 nsew
rlabel metal5 s -8726 624296 592650 624936 6 vssd1
port 538 nsew
rlabel metal5 s -8726 607976 592650 608616 6 vssd1
port 538 nsew
rlabel metal5 s -8726 591656 592650 592296 6 vssd1
port 538 nsew
rlabel metal5 s -8726 575336 592650 575976 6 vssd1
port 538 nsew
rlabel metal5 s -8726 559016 592650 559656 6 vssd1
port 538 nsew
rlabel metal5 s -8726 542696 592650 543336 6 vssd1
port 538 nsew
rlabel metal5 s -8726 526376 592650 527016 6 vssd1
port 538 nsew
rlabel metal5 s -8726 510056 592650 510696 6 vssd1
port 538 nsew
rlabel metal5 s -8726 493736 592650 494376 6 vssd1
port 538 nsew
rlabel metal5 s -8726 477416 592650 478056 6 vssd1
port 538 nsew
rlabel metal5 s -8726 461096 592650 461736 6 vssd1
port 538 nsew
rlabel metal5 s -8726 444776 592650 445416 6 vssd1
port 538 nsew
rlabel metal5 s -8726 428456 592650 429096 6 vssd1
port 538 nsew
rlabel metal5 s -8726 412136 592650 412776 6 vssd1
port 538 nsew
rlabel metal5 s -8726 395816 592650 396456 6 vssd1
port 538 nsew
rlabel metal5 s -8726 379496 592650 380136 6 vssd1
port 538 nsew
rlabel metal5 s -8726 363176 592650 363816 6 vssd1
port 538 nsew
rlabel metal5 s -8726 346856 592650 347496 6 vssd1
port 538 nsew
rlabel metal5 s -8726 330536 592650 331176 6 vssd1
port 538 nsew
rlabel metal5 s -8726 314216 592650 314856 6 vssd1
port 538 nsew
rlabel metal5 s -8726 297896 592650 298536 6 vssd1
port 538 nsew
rlabel metal5 s -8726 281576 592650 282216 6 vssd1
port 538 nsew
rlabel metal5 s -8726 265256 592650 265896 6 vssd1
port 538 nsew
rlabel metal5 s -8726 248936 592650 249576 6 vssd1
port 538 nsew
rlabel metal5 s -8726 232616 592650 233256 6 vssd1
port 538 nsew
rlabel metal5 s -8726 216296 592650 216936 6 vssd1
port 538 nsew
rlabel metal5 s -8726 199976 592650 200616 6 vssd1
port 538 nsew
rlabel metal5 s -8726 183656 592650 184296 6 vssd1
port 538 nsew
rlabel metal5 s -8726 167336 592650 167976 6 vssd1
port 538 nsew
rlabel metal5 s -8726 151016 592650 151656 6 vssd1
port 538 nsew
rlabel metal5 s -8726 134696 592650 135336 6 vssd1
port 538 nsew
rlabel metal5 s -8726 118376 592650 119016 6 vssd1
port 538 nsew
rlabel metal5 s -8726 102056 592650 102696 6 vssd1
port 538 nsew
rlabel metal5 s -8726 85736 592650 86376 6 vssd1
port 538 nsew
rlabel metal5 s -8726 69416 592650 70056 6 vssd1
port 538 nsew
rlabel metal5 s -8726 53096 592650 53736 6 vssd1
port 538 nsew
rlabel metal5 s -8726 36776 592650 37416 6 vssd1
port 538 nsew
rlabel metal5 s -8726 20456 592650 21096 6 vssd1
port 538 nsew
rlabel metal5 s -8726 4136 592650 4776 6 vssd1
port 538 nsew
rlabel metal4 s 574264 -7654 574904 711590 6 vssd1
port 538 nsew
rlabel metal4 s 557944 -7654 558584 711590 6 vssd1
port 538 nsew
rlabel metal4 s 541624 -7654 542264 711590 6 vssd1
port 538 nsew
rlabel metal4 s 525304 -7654 525944 711590 6 vssd1
port 538 nsew
rlabel metal4 s 508984 -7654 509624 711590 6 vssd1
port 538 nsew
rlabel metal4 s 492664 -7654 493304 711590 6 vssd1
port 538 nsew
rlabel metal4 s 476344 -7654 476984 711590 6 vssd1
port 538 nsew
rlabel metal4 s 460024 -7654 460664 711590 6 vssd1
port 538 nsew
rlabel metal4 s 443704 -7654 444344 711590 6 vssd1
port 538 nsew
rlabel metal4 s 427384 -7654 428024 711590 6 vssd1
port 538 nsew
rlabel metal4 s 411064 -7654 411704 711590 6 vssd1
port 538 nsew
rlabel metal4 s 394744 -7654 395384 711590 6 vssd1
port 538 nsew
rlabel metal4 s 378424 -7654 379064 711590 6 vssd1
port 538 nsew
rlabel metal4 s 362104 -7654 362744 711590 6 vssd1
port 538 nsew
rlabel metal4 s 345784 -7654 346424 711590 6 vssd1
port 538 nsew
rlabel metal4 s 329464 -7654 330104 711590 6 vssd1
port 538 nsew
rlabel metal4 s 313144 -7654 313784 711590 6 vssd1
port 538 nsew
rlabel metal4 s 296824 -7654 297464 711590 6 vssd1
port 538 nsew
rlabel metal4 s 280504 -7654 281144 711590 6 vssd1
port 538 nsew
rlabel metal4 s 264184 -7654 264824 711590 6 vssd1
port 538 nsew
rlabel metal4 s 247864 -7654 248504 711590 6 vssd1
port 538 nsew
rlabel metal4 s 231544 -7654 232184 711590 6 vssd1
port 538 nsew
rlabel metal4 s 215224 -7654 215864 711590 6 vssd1
port 538 nsew
rlabel metal4 s 198904 -7654 199544 711590 6 vssd1
port 538 nsew
rlabel metal4 s 182584 -7654 183224 711590 6 vssd1
port 538 nsew
rlabel metal4 s 166264 -7654 166904 711590 6 vssd1
port 538 nsew
rlabel metal4 s 149944 151257 150584 711590 6 vssd1
port 538 nsew
rlabel metal4 s 149944 -7654 150584 4575 8 vssd1
port 538 nsew
rlabel metal4 s 133624 151257 134264 711590 6 vssd1
port 538 nsew
rlabel metal4 s 133624 -7654 134264 4575 8 vssd1
port 538 nsew
rlabel metal4 s 117304 151257 117944 711590 6 vssd1
port 538 nsew
rlabel metal4 s 117304 -7654 117944 4575 8 vssd1
port 538 nsew
rlabel metal4 s 100984 151257 101624 711590 6 vssd1
port 538 nsew
rlabel metal4 s 100984 -7654 101624 4575 8 vssd1
port 538 nsew
rlabel metal4 s 84664 151257 85304 711590 6 vssd1
port 538 nsew
rlabel metal4 s 84664 -7654 85304 4575 8 vssd1
port 538 nsew
rlabel metal4 s 68344 151257 68984 711590 6 vssd1
port 538 nsew
rlabel metal4 s 68344 -7654 68984 4575 8 vssd1
port 538 nsew
rlabel metal4 s 52024 151257 52664 711590 6 vssd1
port 538 nsew
rlabel metal4 s 52024 -7654 52664 4575 8 vssd1
port 538 nsew
rlabel metal4 s 35704 151257 36344 711590 6 vssd1
port 538 nsew
rlabel metal4 s 35704 -7654 36344 4575 8 vssd1
port 538 nsew
rlabel metal4 s 19384 151257 20024 711590 6 vssd1
port 538 nsew
rlabel metal4 s 19384 -7654 20024 4575 8 vssd1
port 538 nsew
rlabel metal4 s 3064 -7654 3704 711590 6 vssd1
port 538 nsew
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew
rlabel metal5 s -8726 692136 592650 692776 6 vssd2
port 539 nsew
rlabel metal5 s -8726 675816 592650 676456 6 vssd2
port 539 nsew
rlabel metal5 s -8726 659496 592650 660136 6 vssd2
port 539 nsew
rlabel metal5 s -8726 643176 592650 643816 6 vssd2
port 539 nsew
rlabel metal5 s -8726 626856 592650 627496 6 vssd2
port 539 nsew
rlabel metal5 s -8726 610536 592650 611176 6 vssd2
port 539 nsew
rlabel metal5 s -8726 594216 592650 594856 6 vssd2
port 539 nsew
rlabel metal5 s -8726 577896 592650 578536 6 vssd2
port 539 nsew
rlabel metal5 s -8726 561576 592650 562216 6 vssd2
port 539 nsew
rlabel metal5 s -8726 545256 592650 545896 6 vssd2
port 539 nsew
rlabel metal5 s -8726 528936 592650 529576 6 vssd2
port 539 nsew
rlabel metal5 s -8726 512616 592650 513256 6 vssd2
port 539 nsew
rlabel metal5 s -8726 496296 592650 496936 6 vssd2
port 539 nsew
rlabel metal5 s -8726 479976 592650 480616 6 vssd2
port 539 nsew
rlabel metal5 s -8726 463656 592650 464296 6 vssd2
port 539 nsew
rlabel metal5 s -8726 447336 592650 447976 6 vssd2
port 539 nsew
rlabel metal5 s -8726 431016 592650 431656 6 vssd2
port 539 nsew
rlabel metal5 s -8726 414696 592650 415336 6 vssd2
port 539 nsew
rlabel metal5 s -8726 398376 592650 399016 6 vssd2
port 539 nsew
rlabel metal5 s -8726 382056 592650 382696 6 vssd2
port 539 nsew
rlabel metal5 s -8726 365736 592650 366376 6 vssd2
port 539 nsew
rlabel metal5 s -8726 349416 592650 350056 6 vssd2
port 539 nsew
rlabel metal5 s -8726 333096 592650 333736 6 vssd2
port 539 nsew
rlabel metal5 s -8726 316776 592650 317416 6 vssd2
port 539 nsew
rlabel metal5 s -8726 300456 592650 301096 6 vssd2
port 539 nsew
rlabel metal5 s -8726 284136 592650 284776 6 vssd2
port 539 nsew
rlabel metal5 s -8726 267816 592650 268456 6 vssd2
port 539 nsew
rlabel metal5 s -8726 251496 592650 252136 6 vssd2
port 539 nsew
rlabel metal5 s -8726 235176 592650 235816 6 vssd2
port 539 nsew
rlabel metal5 s -8726 218856 592650 219496 6 vssd2
port 539 nsew
rlabel metal5 s -8726 202536 592650 203176 6 vssd2
port 539 nsew
rlabel metal5 s -8726 186216 592650 186856 6 vssd2
port 539 nsew
rlabel metal5 s -8726 169896 592650 170536 6 vssd2
port 539 nsew
rlabel metal5 s -8726 153576 592650 154216 6 vssd2
port 539 nsew
rlabel metal5 s -8726 137256 592650 137896 6 vssd2
port 539 nsew
rlabel metal5 s -8726 120936 592650 121576 6 vssd2
port 539 nsew
rlabel metal5 s -8726 104616 592650 105256 6 vssd2
port 539 nsew
rlabel metal5 s -8726 88296 592650 88936 6 vssd2
port 539 nsew
rlabel metal5 s -8726 71976 592650 72616 6 vssd2
port 539 nsew
rlabel metal5 s -8726 55656 592650 56296 6 vssd2
port 539 nsew
rlabel metal5 s -8726 39336 592650 39976 6 vssd2
port 539 nsew
rlabel metal5 s -8726 23016 592650 23656 6 vssd2
port 539 nsew
rlabel metal5 s -8726 6696 592650 7336 6 vssd2
port 539 nsew
rlabel metal4 s 576824 -7654 577464 711590 6 vssd2
port 539 nsew
rlabel metal4 s 560504 -7654 561144 711590 6 vssd2
port 539 nsew
rlabel metal4 s 544184 -7654 544824 711590 6 vssd2
port 539 nsew
rlabel metal4 s 527864 -7654 528504 711590 6 vssd2
port 539 nsew
rlabel metal4 s 511544 -7654 512184 711590 6 vssd2
port 539 nsew
rlabel metal4 s 495224 -7654 495864 711590 6 vssd2
port 539 nsew
rlabel metal4 s 478904 -7654 479544 711590 6 vssd2
port 539 nsew
rlabel metal4 s 462584 -7654 463224 711590 6 vssd2
port 539 nsew
rlabel metal4 s 446264 -7654 446904 711590 6 vssd2
port 539 nsew
rlabel metal4 s 429944 -7654 430584 711590 6 vssd2
port 539 nsew
rlabel metal4 s 413624 -7654 414264 711590 6 vssd2
port 539 nsew
rlabel metal4 s 397304 -7654 397944 711590 6 vssd2
port 539 nsew
rlabel metal4 s 380984 -7654 381624 711590 6 vssd2
port 539 nsew
rlabel metal4 s 364664 -7654 365304 711590 6 vssd2
port 539 nsew
rlabel metal4 s 348344 -7654 348984 711590 6 vssd2
port 539 nsew
rlabel metal4 s 332024 -7654 332664 711590 6 vssd2
port 539 nsew
rlabel metal4 s 315704 -7654 316344 711590 6 vssd2
port 539 nsew
rlabel metal4 s 299384 -7654 300024 711590 6 vssd2
port 539 nsew
rlabel metal4 s 283064 -7654 283704 711590 6 vssd2
port 539 nsew
rlabel metal4 s 266744 -7654 267384 711590 6 vssd2
port 539 nsew
rlabel metal4 s 250424 -7654 251064 711590 6 vssd2
port 539 nsew
rlabel metal4 s 234104 -7654 234744 711590 6 vssd2
port 539 nsew
rlabel metal4 s 217784 -7654 218424 711590 6 vssd2
port 539 nsew
rlabel metal4 s 201464 -7654 202104 711590 6 vssd2
port 539 nsew
rlabel metal4 s 185144 -7654 185784 711590 6 vssd2
port 539 nsew
rlabel metal4 s 168824 -7654 169464 711590 6 vssd2
port 539 nsew
rlabel metal4 s 152504 161888 153144 711590 6 vssd2
port 539 nsew
rlabel metal4 s 136184 161888 136824 711590 6 vssd2
port 539 nsew
rlabel metal4 s 119864 161888 120504 711590 6 vssd2
port 539 nsew
rlabel metal4 s 103544 161888 104184 711590 6 vssd2
port 539 nsew
rlabel metal4 s 87224 161888 87864 711590 6 vssd2
port 539 nsew
rlabel metal4 s 70904 161888 71544 711590 6 vssd2
port 539 nsew
rlabel metal4 s 54584 161888 55224 711590 6 vssd2
port 539 nsew
rlabel metal4 s 38264 161888 38904 711590 6 vssd2
port 539 nsew
rlabel metal4 s 21944 161888 22584 711590 6 vssd2
port 539 nsew
rlabel metal4 s 5624 161888 6264 711590 6 vssd2
port 539 nsew
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 85458310
string GDS_FILE /home/hosni/AES/caravel_aes_example/openlane/user_project_wrapper/runs/23_06_05_14_48/results/signoff/user_project_wrapper.magic.gds
string GDS_START 81748960
<< end >>

