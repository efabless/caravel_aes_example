VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    PORT
      LAYER met5 ;
        RECT -43.630 3441.480 2963.250 3444.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3359.880 2963.250 3363.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3278.280 2963.250 3281.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3196.680 2963.250 3199.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3115.080 2963.250 3118.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3033.480 2963.250 3036.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2951.880 2963.250 2955.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2870.280 2963.250 2873.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2788.680 2963.250 2791.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2707.080 2963.250 2710.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2625.480 2963.250 2628.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2543.880 2963.250 2547.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2462.280 2963.250 2465.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2380.680 2963.250 2383.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2299.080 2963.250 2302.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2217.480 2963.250 2220.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2135.880 2963.250 2139.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2054.280 2963.250 2057.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1972.680 2963.250 1975.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1891.080 2963.250 1894.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1809.480 2963.250 1812.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1727.880 2963.250 1731.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1646.280 2963.250 1649.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1564.680 2963.250 1567.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1483.080 2963.250 1486.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1401.480 2963.250 1404.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1319.880 2963.250 1323.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1238.280 2963.250 1241.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1156.680 2963.250 1159.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1075.080 2963.250 1078.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 993.480 2963.250 996.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 911.880 2963.250 915.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 830.280 2963.250 833.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 748.680 2963.250 751.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 667.080 2963.250 670.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 585.480 2963.250 588.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 503.880 2963.250 507.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 422.280 2963.250 425.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 340.680 2963.250 343.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 259.080 2963.250 262.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 177.480 2963.250 180.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 95.880 2963.250 99.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 14.280 2963.250 17.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 2864.920 -38.270 2868.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2783.320 -38.270 2786.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2701.720 -38.270 2704.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2620.120 -38.270 2623.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2538.520 -38.270 2541.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2456.920 -38.270 2460.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.320 -38.270 2378.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2293.720 -38.270 2296.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2212.120 -38.270 2215.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2130.520 -38.270 2133.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2048.920 -38.270 2052.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1967.320 -38.270 1970.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1885.720 -38.270 1888.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.120 -38.270 1807.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1722.520 -38.270 1725.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1640.920 -38.270 1644.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1559.320 -38.270 1562.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1477.720 -38.270 1480.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.120 -38.270 1399.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1314.520 -38.270 1317.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1232.920 -38.270 1236.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1151.320 -38.270 1154.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1069.720 -38.270 1072.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 988.120 -38.270 991.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.520 -38.270 909.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 824.920 764.445 828.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 824.920 -38.270 828.120 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.320 764.445 746.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.320 -38.270 746.520 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.720 764.445 664.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.720 -38.270 664.920 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 580.120 764.445 583.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 580.120 -38.270 583.320 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.520 764.445 501.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.520 -38.270 501.720 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.920 764.445 420.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.920 -38.270 420.120 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.320 764.445 338.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.320 -38.270 338.520 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 253.720 764.445 256.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 253.720 -38.270 256.920 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 172.120 764.445 175.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 172.120 -38.270 175.320 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.520 764.445 93.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.520 -38.270 93.720 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.920 -38.270 12.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
  END vccd1
  PIN vccd2
    PORT
      LAYER met5 ;
        RECT -43.630 3454.280 2963.250 3457.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3372.680 2963.250 3375.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3291.080 2963.250 3294.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3209.480 2963.250 3212.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3127.880 2963.250 3131.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3046.280 2963.250 3049.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2964.680 2963.250 2967.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2883.080 2963.250 2886.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2801.480 2963.250 2804.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2719.880 2963.250 2723.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2638.280 2963.250 2641.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2556.680 2963.250 2559.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2475.080 2963.250 2478.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2393.480 2963.250 2396.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2311.880 2963.250 2315.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.280 2963.250 2233.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2148.680 2963.250 2151.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2067.080 2963.250 2070.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1985.480 2963.250 1988.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1903.880 2963.250 1907.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1822.280 2963.250 1825.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1740.680 2963.250 1743.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1659.080 2963.250 1662.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1577.480 2963.250 1580.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1495.880 2963.250 1499.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1414.280 2963.250 1417.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1332.680 2963.250 1335.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1251.080 2963.250 1254.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1169.480 2963.250 1172.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1087.880 2963.250 1091.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1006.280 2963.250 1009.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 924.680 2963.250 927.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 843.080 2963.250 846.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 761.480 2963.250 764.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 679.880 2963.250 683.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 598.280 2963.250 601.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 516.680 2963.250 519.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 435.080 2963.250 438.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 353.480 2963.250 356.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 271.880 2963.250 275.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 190.280 2963.250 193.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 108.680 2963.250 111.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 27.080 2963.250 30.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2877.720 -38.270 2880.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2796.120 -38.270 2799.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2714.520 -38.270 2717.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.920 -38.270 2636.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2551.320 -38.270 2554.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2469.720 -38.270 2472.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2388.120 -38.270 2391.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2306.520 -38.270 2309.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.920 -38.270 2228.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2143.320 -38.270 2146.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.720 -38.270 2064.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.120 -38.270 1983.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.520 -38.270 1901.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1816.920 -38.270 1820.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.320 -38.270 1738.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1653.720 -38.270 1656.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1572.120 -38.270 1575.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1490.520 -38.270 1493.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.920 -38.270 1412.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1327.320 -38.270 1330.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1245.720 -38.270 1248.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.120 -38.270 1167.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1082.520 -38.270 1085.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1000.920 -38.270 1004.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 919.320 -38.270 922.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.720 -38.270 840.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.120 764.445 759.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.520 764.445 677.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 592.920 764.445 596.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 511.320 764.445 514.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 429.720 764.445 432.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 348.120 764.445 351.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 266.520 764.445 269.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.920 764.445 188.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.320 764.445 106.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.720 764.445 24.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
  END vccd2
  PIN vdda1
    PORT
      LAYER met5 ;
        RECT -43.630 3467.080 2963.250 3470.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3385.480 2963.250 3388.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3303.880 2963.250 3307.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3222.280 2963.250 3225.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3140.680 2963.250 3143.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3059.080 2963.250 3062.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2977.480 2963.250 2980.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2895.880 2963.250 2899.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2814.280 2963.250 2817.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2732.680 2963.250 2735.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2651.080 2963.250 2654.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2569.480 2963.250 2572.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2487.880 2963.250 2491.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2406.280 2963.250 2409.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2324.680 2963.250 2327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2243.080 2963.250 2246.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2161.480 2963.250 2164.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2079.880 2963.250 2083.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1998.280 2963.250 2001.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1916.680 2963.250 1919.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1835.080 2963.250 1838.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1753.480 2963.250 1756.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1671.880 2963.250 1675.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1590.280 2963.250 1593.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1508.680 2963.250 1511.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1427.080 2963.250 1430.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1345.480 2963.250 1348.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1263.880 2963.250 1267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1182.280 2963.250 1185.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1100.680 2963.250 1103.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1019.080 2963.250 1022.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 937.480 2963.250 940.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 855.880 2963.250 859.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 774.280 2963.250 777.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 692.680 2963.250 695.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 611.080 2963.250 614.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 529.480 2963.250 532.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 447.880 2963.250 451.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 366.280 2963.250 369.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 284.680 2963.250 287.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 203.080 2963.250 206.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 121.480 2963.250 124.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 39.880 2963.250 43.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2890.520 -38.270 2893.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.920 -38.270 2812.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.320 -38.270 2730.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2645.720 -38.270 2648.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2564.120 -38.270 2567.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2482.520 -38.270 2485.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2400.920 -38.270 2404.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2319.320 -38.270 2322.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2237.720 -38.270 2240.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.120 -38.270 2159.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.520 -38.270 2077.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1992.920 -38.270 1996.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.320 -38.270 1914.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.720 -38.270 1832.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1748.120 -38.270 1751.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.520 -38.270 1669.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.920 -38.270 1588.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1503.320 -38.270 1506.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.720 -38.270 1424.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1340.120 -38.270 1343.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.520 -38.270 1261.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1176.920 -38.270 1180.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.320 -38.270 1098.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.720 -38.270 1016.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.120 -38.270 935.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 850.520 -38.270 853.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 768.920 764.445 772.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 687.320 764.445 690.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.720 764.445 608.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.120 764.445 527.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 442.520 764.445 445.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 360.920 764.445 364.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.320 764.445 282.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.720 764.445 200.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.120 764.445 119.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.520 764.445 37.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
  END vdda1
  PIN vdda2
    PORT
      LAYER met5 ;
        RECT -43.630 3479.880 2963.250 3483.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3398.280 2963.250 3401.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3316.680 2963.250 3319.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3235.080 2963.250 3238.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3153.480 2963.250 3156.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3071.880 2963.250 3075.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2990.280 2963.250 2993.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2908.680 2963.250 2911.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2827.080 2963.250 2830.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2745.480 2963.250 2748.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2663.880 2963.250 2667.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2582.280 2963.250 2585.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2500.680 2963.250 2503.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2419.080 2963.250 2422.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2337.480 2963.250 2340.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2255.880 2963.250 2259.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2174.280 2963.250 2177.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2092.680 2963.250 2095.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2011.080 2963.250 2014.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1929.480 2963.250 1932.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1847.880 2963.250 1851.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1766.280 2963.250 1769.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1684.680 2963.250 1687.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1603.080 2963.250 1606.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1521.480 2963.250 1524.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1439.880 2963.250 1443.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1358.280 2963.250 1361.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1276.680 2963.250 1279.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1195.080 2963.250 1198.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1113.480 2963.250 1116.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1031.880 2963.250 1035.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 950.280 2963.250 953.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 868.680 2963.250 871.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 787.080 2963.250 790.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 705.480 2963.250 708.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 623.880 2963.250 627.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 542.280 2963.250 545.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 460.680 2963.250 463.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 379.080 2963.250 382.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 297.480 2963.250 300.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 215.880 2963.250 219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 134.280 2963.250 137.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 52.680 2963.250 55.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2903.320 -38.270 2906.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2821.720 -38.270 2824.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2740.120 -38.270 2743.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.520 -38.270 2661.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2576.920 -38.270 2580.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2495.320 -38.270 2498.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2413.720 -38.270 2416.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.120 -38.270 2335.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2250.520 -38.270 2253.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.920 -38.270 2172.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2087.320 -38.270 2090.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2005.720 -38.270 2008.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1924.120 -38.270 1927.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1842.520 -38.270 1845.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1760.920 -38.270 1764.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1679.320 -38.270 1682.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1597.720 -38.270 1600.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.120 -38.270 1519.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.520 -38.270 1437.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1352.920 -38.270 1356.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.320 -38.270 1274.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1189.720 -38.270 1192.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.120 -38.270 1111.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.520 -38.270 1029.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 944.920 -38.270 948.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.320 -38.270 866.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 781.720 764.445 784.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.120 764.445 703.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 618.520 764.445 621.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 536.920 764.445 540.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 455.320 764.445 458.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 373.720 764.445 376.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 292.120 764.445 295.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 210.520 764.445 213.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.920 764.445 132.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.320 764.445 50.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
  END vdda2
  PIN vssa1
    PORT
      LAYER met5 ;
        RECT -43.630 3473.480 2963.250 3476.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3391.880 2963.250 3395.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.280 2963.250 3313.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3228.680 2963.250 3231.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3147.080 2963.250 3150.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3065.480 2963.250 3068.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2983.880 2963.250 2987.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2902.280 2963.250 2905.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2820.680 2963.250 2823.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2739.080 2963.250 2742.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2657.480 2963.250 2660.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2575.880 2963.250 2579.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2494.280 2963.250 2497.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2412.680 2963.250 2415.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2331.080 2963.250 2334.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2249.480 2963.250 2252.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2167.880 2963.250 2171.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2086.280 2963.250 2089.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2004.680 2963.250 2007.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1923.080 2963.250 1926.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1841.480 2963.250 1844.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1759.880 2963.250 1763.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1678.280 2963.250 1681.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1596.680 2963.250 1599.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1515.080 2963.250 1518.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1433.480 2963.250 1436.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1351.880 2963.250 1355.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1270.280 2963.250 1273.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1188.680 2963.250 1191.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1107.080 2963.250 1110.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1025.480 2963.250 1028.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 943.880 2963.250 947.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 862.280 2963.250 865.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 780.680 2963.250 783.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 699.080 2963.250 702.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 617.480 2963.250 620.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 535.880 2963.250 539.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 454.280 2963.250 457.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 372.680 2963.250 375.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 291.080 2963.250 294.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 209.480 2963.250 212.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 127.880 2963.250 131.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 46.280 2963.250 49.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 2896.920 -38.270 2900.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2815.320 -38.270 2818.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2733.720 -38.270 2736.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2652.120 -38.270 2655.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2570.520 -38.270 2573.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2488.920 -38.270 2492.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2407.320 -38.270 2410.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.720 -38.270 2328.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2244.120 -38.270 2247.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2162.520 -38.270 2165.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2080.920 -38.270 2084.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1999.320 -38.270 2002.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.720 -38.270 1920.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1836.120 -38.270 1839.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1754.520 -38.270 1757.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1672.920 -38.270 1676.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1591.320 -38.270 1594.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1509.720 -38.270 1512.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1428.120 -38.270 1431.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.520 -38.270 1349.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.920 -38.270 1268.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1183.320 -38.270 1186.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1101.720 -38.270 1104.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1020.120 -38.270 1023.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 938.520 -38.270 941.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.920 -38.270 860.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.320 764.445 778.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.720 764.445 696.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 612.120 764.445 615.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 530.520 764.445 533.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.920 764.445 452.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 367.320 764.445 370.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 285.720 764.445 288.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.120 764.445 207.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.520 764.445 125.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.920 764.445 44.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
  END vssa1
  PIN vssa2
    PORT
      LAYER met5 ;
        RECT -43.630 3486.280 2963.250 3489.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3404.680 2963.250 3407.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3323.080 2963.250 3326.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3241.480 2963.250 3244.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3159.880 2963.250 3163.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3078.280 2963.250 3081.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2996.680 2963.250 2999.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2915.080 2963.250 2918.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2833.480 2963.250 2836.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2751.880 2963.250 2755.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2670.280 2963.250 2673.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2588.680 2963.250 2591.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2507.080 2963.250 2510.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2425.480 2963.250 2428.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2343.880 2963.250 2347.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2262.280 2963.250 2265.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2180.680 2963.250 2183.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2099.080 2963.250 2102.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2017.480 2963.250 2020.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1935.880 2963.250 1939.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1854.280 2963.250 1857.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1772.680 2963.250 1775.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1691.080 2963.250 1694.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1609.480 2963.250 1612.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1527.880 2963.250 1531.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1446.280 2963.250 1449.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1364.680 2963.250 1367.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1283.080 2963.250 1286.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1201.480 2963.250 1204.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1119.880 2963.250 1123.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1038.280 2963.250 1041.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 956.680 2963.250 959.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 875.080 2963.250 878.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 793.480 2963.250 796.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 711.880 2963.250 715.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 630.280 2963.250 633.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 548.680 2963.250 551.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 467.080 2963.250 470.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 385.480 2963.250 388.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 303.880 2963.250 307.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 222.280 2963.250 225.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 140.680 2963.250 143.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 59.080 2963.250 62.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2909.720 -38.270 2912.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2828.120 -38.270 2831.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.520 -38.270 2749.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.920 -38.270 2668.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2583.320 -38.270 2586.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2501.720 -38.270 2504.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2420.120 -38.270 2423.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2338.520 -38.270 2341.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2256.920 -38.270 2260.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.320 -38.270 2178.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2093.720 -38.270 2096.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2012.120 -38.270 2015.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1930.520 -38.270 1933.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1848.920 -38.270 1852.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1767.320 -38.270 1770.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1685.720 -38.270 1688.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.120 -38.270 1607.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1522.520 -38.270 1525.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1440.920 -38.270 1444.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1359.320 -38.270 1362.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1277.720 -38.270 1280.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1196.120 -38.270 1199.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.520 -38.270 1117.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.920 -38.270 1036.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.320 -38.270 954.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 869.720 -38.270 872.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 788.120 764.445 791.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.520 764.445 709.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.920 764.445 628.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 543.320 764.445 546.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 764.445 464.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 380.120 764.445 383.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 298.520 764.445 301.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.920 764.445 220.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.320 764.445 138.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.720 764.445 56.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
  END vssa2
  PIN vssd1
    PORT
      LAYER met5 ;
        RECT -43.630 3447.880 2963.250 3451.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3366.280 2963.250 3369.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3284.680 2963.250 3287.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3203.080 2963.250 3206.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3121.480 2963.250 3124.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3039.880 2963.250 3043.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2958.280 2963.250 2961.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2876.680 2963.250 2879.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2795.080 2963.250 2798.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2713.480 2963.250 2716.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2631.880 2963.250 2635.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2550.280 2963.250 2553.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2468.680 2963.250 2471.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2387.080 2963.250 2390.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2305.480 2963.250 2308.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2223.880 2963.250 2227.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2142.280 2963.250 2145.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2060.680 2963.250 2063.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1979.080 2963.250 1982.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1897.480 2963.250 1900.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1815.880 2963.250 1819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1734.280 2963.250 1737.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1652.680 2963.250 1655.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1571.080 2963.250 1574.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1489.480 2963.250 1492.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1407.880 2963.250 1411.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1326.280 2963.250 1329.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1244.680 2963.250 1247.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1163.080 2963.250 1166.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1081.480 2963.250 1084.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 999.880 2963.250 1003.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 918.280 2963.250 921.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 836.680 2963.250 839.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 755.080 2963.250 758.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 673.480 2963.250 676.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 591.880 2963.250 595.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 510.280 2963.250 513.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 428.680 2963.250 431.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 347.080 2963.250 350.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 265.480 2963.250 268.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 183.880 2963.250 187.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 102.280 2963.250 105.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 20.680 2963.250 23.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2871.320 -38.270 2874.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2789.720 -38.270 2792.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.120 -38.270 2711.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2626.520 -38.270 2629.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2544.920 -38.270 2548.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2463.320 -38.270 2466.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2381.720 -38.270 2384.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2300.120 -38.270 2303.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2218.520 -38.270 2221.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2136.920 -38.270 2140.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.320 -38.270 2058.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1973.720 -38.270 1976.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1892.120 -38.270 1895.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1810.520 -38.270 1813.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.920 -38.270 1732.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.320 -38.270 1650.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1565.720 -38.270 1568.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1484.120 -38.270 1487.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1402.520 -38.270 1405.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1320.920 -38.270 1324.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1239.320 -38.270 1242.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1157.720 -38.270 1160.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1076.120 -38.270 1079.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 994.520 -38.270 997.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 912.920 -38.270 916.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.320 -38.270 834.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 749.720 764.445 752.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 749.720 -38.270 752.920 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.120 764.445 671.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.120 -38.270 671.320 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.520 764.445 589.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.520 -38.270 589.720 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.920 764.445 508.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.920 -38.270 508.120 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.320 764.445 426.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.320 -38.270 426.520 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.720 764.445 344.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.720 -38.270 344.920 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 260.120 764.445 263.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 260.120 -38.270 263.320 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 178.520 764.445 181.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 178.520 -38.270 181.720 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.920 764.445 100.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.920 -38.270 100.120 24.915 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.320 -38.270 18.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
  END vssd1
  PIN vssd2
    PORT
      LAYER met5 ;
        RECT -43.630 3460.680 2963.250 3463.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3379.080 2963.250 3382.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3297.480 2963.250 3300.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3215.880 2963.250 3219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3134.280 2963.250 3137.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3052.680 2963.250 3055.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2971.080 2963.250 2974.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2889.480 2963.250 2892.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2807.880 2963.250 2811.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2726.280 2963.250 2729.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2644.680 2963.250 2647.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2563.080 2963.250 2566.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2481.480 2963.250 2484.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2399.880 2963.250 2403.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2318.280 2963.250 2321.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2236.680 2963.250 2239.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2155.080 2963.250 2158.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2073.480 2963.250 2076.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1991.880 2963.250 1995.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1910.280 2963.250 1913.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1828.680 2963.250 1831.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1747.080 2963.250 1750.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1665.480 2963.250 1668.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1583.880 2963.250 1587.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1502.280 2963.250 1505.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.680 2963.250 1423.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1339.080 2963.250 1342.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1257.480 2963.250 1260.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1175.880 2963.250 1179.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1094.280 2963.250 1097.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1012.680 2963.250 1015.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 931.080 2963.250 934.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 849.480 2963.250 852.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 767.880 2963.250 771.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 686.280 2963.250 689.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 604.680 2963.250 607.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 523.080 2963.250 526.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 441.480 2963.250 444.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 359.880 2963.250 363.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 278.280 2963.250 281.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 196.680 2963.250 199.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 115.080 2963.250 118.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 33.480 2963.250 36.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2884.120 -38.270 2887.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2802.520 -38.270 2805.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2720.920 -38.270 2724.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2639.320 -38.270 2642.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2557.720 -38.270 2560.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.120 -38.270 2479.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.520 -38.270 2397.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2312.920 -38.270 2316.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.320 -38.270 2234.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2149.720 -38.270 2152.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2068.120 -38.270 2071.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1986.520 -38.270 1989.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.920 -38.270 1908.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.320 -38.270 1826.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1741.720 -38.270 1744.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1660.120 -38.270 1663.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1578.520 -38.270 1581.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.920 -38.270 1500.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.320 -38.270 1418.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1333.720 -38.270 1336.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1252.120 -38.270 1255.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1170.520 -38.270 1173.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.920 -38.270 1092.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.320 -38.270 1010.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 925.720 -38.270 928.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 844.120 -38.270 847.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 762.520 809.440 765.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 680.920 809.440 684.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.320 809.440 602.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 517.720 809.440 520.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.120 809.440 439.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.520 809.440 357.720 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 272.920 809.440 276.120 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.320 809.440 194.520 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 109.720 809.440 112.920 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.120 809.440 31.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 15.520 30.795 824.200 808.885 ;
      LAYER met1 ;
        RECT 15.520 10.240 826.430 809.040 ;
      LAYER met2 ;
        RECT 2.850 2.680 826.400 808.985 ;
        RECT 3.550 1.630 7.950 2.680 ;
        RECT 9.070 1.630 13.930 2.680 ;
        RECT 15.050 1.630 19.910 2.680 ;
        RECT 21.030 1.630 25.890 2.680 ;
        RECT 27.010 1.630 31.870 2.680 ;
        RECT 32.990 1.630 37.850 2.680 ;
        RECT 38.970 1.630 43.370 2.680 ;
        RECT 44.490 1.630 49.350 2.680 ;
        RECT 50.470 1.630 55.330 2.680 ;
        RECT 56.450 1.630 61.310 2.680 ;
        RECT 62.430 1.630 67.290 2.680 ;
        RECT 68.410 1.630 73.270 2.680 ;
        RECT 74.390 1.630 79.250 2.680 ;
        RECT 80.370 1.630 84.770 2.680 ;
        RECT 85.890 1.630 90.750 2.680 ;
        RECT 91.870 1.630 96.730 2.680 ;
        RECT 97.850 1.630 102.710 2.680 ;
        RECT 103.830 1.630 108.690 2.680 ;
        RECT 109.810 1.630 114.670 2.680 ;
        RECT 115.790 1.630 120.650 2.680 ;
        RECT 121.770 1.630 126.170 2.680 ;
        RECT 127.290 1.630 132.150 2.680 ;
        RECT 133.270 1.630 138.130 2.680 ;
        RECT 139.250 1.630 144.110 2.680 ;
        RECT 145.230 1.630 150.090 2.680 ;
        RECT 151.210 1.630 156.070 2.680 ;
        RECT 157.190 1.630 161.590 2.680 ;
        RECT 162.710 1.630 167.570 2.680 ;
        RECT 168.690 1.630 173.550 2.680 ;
        RECT 174.670 1.630 179.530 2.680 ;
        RECT 180.650 1.630 185.510 2.680 ;
        RECT 186.630 1.630 191.490 2.680 ;
        RECT 192.610 1.630 197.470 2.680 ;
        RECT 198.590 1.630 202.990 2.680 ;
        RECT 204.110 1.630 208.970 2.680 ;
        RECT 210.090 1.630 214.950 2.680 ;
        RECT 216.070 1.630 220.930 2.680 ;
        RECT 222.050 1.630 226.910 2.680 ;
        RECT 228.030 1.630 232.890 2.680 ;
        RECT 234.010 1.630 238.870 2.680 ;
        RECT 239.990 1.630 244.390 2.680 ;
        RECT 245.510 1.630 250.370 2.680 ;
        RECT 251.490 1.630 256.350 2.680 ;
        RECT 257.470 1.630 262.330 2.680 ;
        RECT 263.450 1.630 268.310 2.680 ;
        RECT 269.430 1.630 274.290 2.680 ;
        RECT 275.410 1.630 279.810 2.680 ;
        RECT 280.930 1.630 285.790 2.680 ;
        RECT 286.910 1.630 291.770 2.680 ;
        RECT 292.890 1.630 297.750 2.680 ;
        RECT 298.870 1.630 303.730 2.680 ;
        RECT 304.850 1.630 309.710 2.680 ;
        RECT 310.830 1.630 315.690 2.680 ;
        RECT 316.810 1.630 321.210 2.680 ;
        RECT 322.330 1.630 327.190 2.680 ;
        RECT 328.310 1.630 333.170 2.680 ;
        RECT 334.290 1.630 339.150 2.680 ;
        RECT 340.270 1.630 345.130 2.680 ;
        RECT 346.250 1.630 351.110 2.680 ;
        RECT 352.230 1.630 357.090 2.680 ;
        RECT 358.210 1.630 362.610 2.680 ;
        RECT 363.730 1.630 368.590 2.680 ;
        RECT 369.710 1.630 374.570 2.680 ;
        RECT 375.690 1.630 380.550 2.680 ;
        RECT 381.670 1.630 386.530 2.680 ;
        RECT 387.650 1.630 392.510 2.680 ;
        RECT 393.630 1.630 398.030 2.680 ;
        RECT 399.150 1.630 404.010 2.680 ;
        RECT 405.130 1.630 409.990 2.680 ;
        RECT 411.110 1.630 415.970 2.680 ;
        RECT 417.090 1.630 421.950 2.680 ;
        RECT 423.070 1.630 427.930 2.680 ;
        RECT 429.050 1.630 433.910 2.680 ;
        RECT 435.030 1.630 439.430 2.680 ;
        RECT 440.550 1.630 445.410 2.680 ;
        RECT 446.530 1.630 451.390 2.680 ;
        RECT 452.510 1.630 457.370 2.680 ;
        RECT 458.490 1.630 463.350 2.680 ;
        RECT 464.470 1.630 469.330 2.680 ;
        RECT 470.450 1.630 475.310 2.680 ;
        RECT 476.430 1.630 480.830 2.680 ;
        RECT 481.950 1.630 486.810 2.680 ;
        RECT 487.930 1.630 492.790 2.680 ;
        RECT 493.910 1.630 498.770 2.680 ;
        RECT 499.890 1.630 504.750 2.680 ;
        RECT 505.870 1.630 510.730 2.680 ;
        RECT 511.850 1.630 516.250 2.680 ;
        RECT 517.370 1.630 522.230 2.680 ;
        RECT 523.350 1.630 528.210 2.680 ;
        RECT 529.330 1.630 534.190 2.680 ;
        RECT 535.310 1.630 540.170 2.680 ;
        RECT 541.290 1.630 546.150 2.680 ;
        RECT 547.270 1.630 552.130 2.680 ;
        RECT 553.250 1.630 557.650 2.680 ;
        RECT 558.770 1.630 563.630 2.680 ;
        RECT 564.750 1.630 569.610 2.680 ;
        RECT 570.730 1.630 575.590 2.680 ;
        RECT 576.710 1.630 581.570 2.680 ;
        RECT 582.690 1.630 587.550 2.680 ;
        RECT 588.670 1.630 593.530 2.680 ;
        RECT 594.650 1.630 599.050 2.680 ;
        RECT 600.170 1.630 605.030 2.680 ;
        RECT 606.150 1.630 611.010 2.680 ;
        RECT 612.130 1.630 616.990 2.680 ;
        RECT 618.110 1.630 622.970 2.680 ;
        RECT 624.090 1.630 628.950 2.680 ;
        RECT 630.070 1.630 634.470 2.680 ;
        RECT 635.590 1.630 640.450 2.680 ;
        RECT 641.570 1.630 646.430 2.680 ;
        RECT 647.550 1.630 652.410 2.680 ;
        RECT 653.530 1.630 658.390 2.680 ;
        RECT 659.510 1.630 664.370 2.680 ;
        RECT 665.490 1.630 670.350 2.680 ;
        RECT 671.470 1.630 675.870 2.680 ;
        RECT 676.990 1.630 681.850 2.680 ;
        RECT 682.970 1.630 687.830 2.680 ;
        RECT 688.950 1.630 693.810 2.680 ;
        RECT 694.930 1.630 699.790 2.680 ;
        RECT 700.910 1.630 705.770 2.680 ;
        RECT 706.890 1.630 711.750 2.680 ;
        RECT 712.870 1.630 717.270 2.680 ;
        RECT 718.390 1.630 723.250 2.680 ;
        RECT 724.370 1.630 729.230 2.680 ;
        RECT 730.350 1.630 735.210 2.680 ;
        RECT 736.330 1.630 741.190 2.680 ;
        RECT 742.310 1.630 747.170 2.680 ;
        RECT 748.290 1.630 752.690 2.680 ;
        RECT 753.810 1.630 758.670 2.680 ;
        RECT 759.790 1.630 764.650 2.680 ;
        RECT 765.770 1.630 770.630 2.680 ;
        RECT 771.750 1.630 776.610 2.680 ;
        RECT 777.730 1.630 782.590 2.680 ;
        RECT 783.710 1.630 788.570 2.680 ;
        RECT 789.690 1.630 794.090 2.680 ;
        RECT 795.210 1.630 800.070 2.680 ;
        RECT 801.190 1.630 806.050 2.680 ;
        RECT 807.170 1.630 812.030 2.680 ;
        RECT 813.150 1.630 818.010 2.680 ;
        RECT 819.130 1.630 823.990 2.680 ;
        RECT 825.110 1.630 826.400 2.680 ;
      LAYER met3 ;
        RECT 2.825 8.335 825.975 808.965 ;
      LAYER met4 ;
        RECT 30.240 764.045 34.120 809.040 ;
        RECT 38.120 764.045 40.520 809.040 ;
        RECT 44.520 764.045 46.920 809.040 ;
        RECT 50.920 764.045 53.320 809.040 ;
        RECT 57.320 764.045 90.120 809.040 ;
        RECT 94.120 764.045 96.520 809.040 ;
        RECT 100.520 764.045 102.920 809.040 ;
        RECT 106.920 764.045 115.720 809.040 ;
        RECT 119.720 764.045 122.120 809.040 ;
        RECT 126.120 764.045 128.520 809.040 ;
        RECT 132.520 764.045 134.920 809.040 ;
        RECT 138.920 764.045 171.720 809.040 ;
        RECT 175.720 764.045 178.120 809.040 ;
        RECT 182.120 764.045 184.520 809.040 ;
        RECT 188.520 764.045 197.320 809.040 ;
        RECT 201.320 764.045 203.720 809.040 ;
        RECT 207.720 764.045 210.120 809.040 ;
        RECT 214.120 764.045 216.520 809.040 ;
        RECT 220.520 764.045 253.320 809.040 ;
        RECT 257.320 764.045 259.720 809.040 ;
        RECT 263.720 764.045 266.120 809.040 ;
        RECT 270.120 764.045 278.920 809.040 ;
        RECT 282.920 764.045 285.320 809.040 ;
        RECT 289.320 764.045 291.720 809.040 ;
        RECT 295.720 764.045 298.120 809.040 ;
        RECT 302.120 764.045 334.920 809.040 ;
        RECT 338.920 764.045 341.320 809.040 ;
        RECT 345.320 764.045 347.720 809.040 ;
        RECT 351.720 764.045 360.520 809.040 ;
        RECT 364.520 764.045 366.920 809.040 ;
        RECT 370.920 764.045 373.320 809.040 ;
        RECT 377.320 764.045 379.720 809.040 ;
        RECT 383.720 764.045 416.520 809.040 ;
        RECT 420.520 764.045 422.920 809.040 ;
        RECT 426.920 764.045 429.320 809.040 ;
        RECT 433.320 764.045 442.120 809.040 ;
        RECT 446.120 764.045 448.520 809.040 ;
        RECT 452.520 764.045 454.920 809.040 ;
        RECT 458.920 764.045 461.320 809.040 ;
        RECT 465.320 764.045 498.120 809.040 ;
        RECT 502.120 764.045 504.520 809.040 ;
        RECT 508.520 764.045 510.920 809.040 ;
        RECT 514.920 764.045 523.720 809.040 ;
        RECT 527.720 764.045 530.120 809.040 ;
        RECT 534.120 764.045 536.520 809.040 ;
        RECT 540.520 764.045 542.920 809.040 ;
        RECT 546.920 764.045 579.720 809.040 ;
        RECT 583.720 764.045 586.120 809.040 ;
        RECT 590.120 764.045 592.520 809.040 ;
        RECT 596.520 764.045 605.320 809.040 ;
        RECT 609.320 764.045 611.720 809.040 ;
        RECT 615.720 764.045 618.120 809.040 ;
        RECT 622.120 764.045 624.520 809.040 ;
        RECT 628.520 764.045 661.320 809.040 ;
        RECT 665.320 764.045 667.720 809.040 ;
        RECT 671.720 764.045 674.120 809.040 ;
        RECT 678.120 764.045 686.920 809.040 ;
        RECT 690.920 764.045 693.320 809.040 ;
        RECT 697.320 764.045 699.720 809.040 ;
        RECT 703.720 764.045 706.120 809.040 ;
        RECT 710.120 764.045 742.920 809.040 ;
        RECT 746.920 764.045 749.320 809.040 ;
        RECT 753.320 764.045 755.720 809.040 ;
        RECT 759.720 764.045 768.520 809.040 ;
        RECT 772.520 764.045 774.920 809.040 ;
        RECT 778.920 764.045 781.320 809.040 ;
        RECT 785.320 764.045 787.720 809.040 ;
        RECT 791.720 764.045 816.545 809.040 ;
        RECT 30.240 25.615 816.545 764.045 ;
  END
END user_project_wrapper
END LIBRARY

