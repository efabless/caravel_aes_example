magic
tech sky130A
magscale 1 2
timestamp 1686145997
<< nwell >>
rect 1066 156933 162878 157499
rect 1066 155845 162878 156411
rect 1066 154757 162878 155323
rect 1066 153669 162878 154235
rect 1066 152581 162878 153147
rect 1066 151493 162878 152059
rect 1066 150405 162878 150971
rect 1066 149317 162878 149883
rect 1066 148229 162878 148795
rect 1066 147141 162878 147707
rect 1066 146053 162878 146619
rect 1066 144965 162878 145531
rect 1066 143877 162878 144443
rect 1066 142789 162878 143355
rect 1066 141701 162878 142267
rect 1066 140613 162878 141179
rect 1066 139525 162878 140091
rect 1066 138437 162878 139003
rect 1066 137349 162878 137915
rect 1066 136261 162878 136827
rect 1066 135173 162878 135739
rect 1066 134085 162878 134651
rect 1066 132997 162878 133563
rect 1066 131909 162878 132475
rect 1066 130821 162878 131387
rect 1066 129733 162878 130299
rect 1066 128645 162878 129211
rect 1066 127557 162878 128123
rect 1066 126469 162878 127035
rect 1066 125381 162878 125947
rect 1066 124293 162878 124859
rect 1066 123205 162878 123771
rect 1066 122117 162878 122683
rect 1066 121029 162878 121595
rect 1066 119941 162878 120507
rect 1066 118853 162878 119419
rect 1066 117765 162878 118331
rect 1066 116677 162878 117243
rect 1066 115589 162878 116155
rect 1066 114501 162878 115067
rect 1066 113413 162878 113979
rect 1066 112325 162878 112891
rect 1066 111237 162878 111803
rect 1066 110149 162878 110715
rect 1066 109061 162878 109627
rect 1066 107973 162878 108539
rect 1066 106885 162878 107451
rect 1066 105797 162878 106363
rect 1066 104709 162878 105275
rect 1066 103621 162878 104187
rect 1066 102533 162878 103099
rect 1066 101445 162878 102011
rect 1066 100357 162878 100923
rect 1066 99269 162878 99835
rect 1066 98181 162878 98747
rect 1066 97093 162878 97659
rect 1066 96005 162878 96571
rect 1066 94917 162878 95483
rect 1066 93829 162878 94395
rect 1066 92741 162878 93307
rect 1066 91653 162878 92219
rect 1066 90565 162878 91131
rect 1066 89477 162878 90043
rect 1066 88389 162878 88955
rect 1066 87301 162878 87867
rect 1066 86213 162878 86779
rect 1066 85125 162878 85691
rect 1066 84037 162878 84603
rect 1066 82949 162878 83515
rect 1066 81861 162878 82427
rect 1066 80773 162878 81339
rect 1066 79685 162878 80251
rect 1066 78597 162878 79163
rect 1066 77509 162878 78075
rect 1066 76421 162878 76987
rect 1066 75333 162878 75899
rect 1066 74245 162878 74811
rect 1066 73157 162878 73723
rect 1066 72069 162878 72635
rect 1066 70981 162878 71547
rect 1066 69893 162878 70459
rect 1066 68805 162878 69371
rect 1066 67717 162878 68283
rect 1066 66629 162878 67195
rect 1066 65541 162878 66107
rect 1066 64453 162878 65019
rect 1066 63365 162878 63931
rect 1066 62277 162878 62843
rect 1066 61189 162878 61755
rect 1066 60101 162878 60667
rect 1066 59013 162878 59579
rect 1066 57925 162878 58491
rect 1066 56837 162878 57403
rect 1066 55749 162878 56315
rect 1066 54661 162878 55227
rect 1066 53573 162878 54139
rect 1066 52485 162878 53051
rect 1066 51397 162878 51963
rect 1066 50309 162878 50875
rect 1066 49221 162878 49787
rect 1066 48133 162878 48699
rect 1066 47045 162878 47611
rect 1066 45957 162878 46523
rect 1066 44869 162878 45435
rect 1066 43781 162878 44347
rect 1066 42693 162878 43259
rect 1066 41605 162878 42171
rect 1066 40517 162878 41083
rect 1066 39429 162878 39995
rect 1066 38341 162878 38907
rect 1066 37253 162878 37819
rect 1066 36165 162878 36731
rect 1066 35077 162878 35643
rect 1066 33989 162878 34555
rect 1066 32901 162878 33467
rect 1066 31813 162878 32379
rect 1066 30725 162878 31291
rect 1066 29637 162878 30203
rect 1066 28549 162878 29115
rect 1066 27461 162878 28027
rect 1066 26373 162878 26939
rect 1066 25285 162878 25851
rect 1066 24197 162878 24763
rect 1066 23109 162878 23675
rect 1066 22021 162878 22587
rect 1066 20933 162878 21499
rect 1066 19845 162878 20411
rect 1066 18757 162878 19323
rect 1066 17669 162878 18235
rect 1066 16581 162878 17147
rect 1066 15493 162878 16059
rect 1066 14405 162878 14971
rect 1066 13317 162878 13883
rect 1066 12229 162878 12795
rect 1066 11141 162878 11707
rect 1066 10053 162878 10619
rect 1066 8965 162878 9531
rect 1066 7877 162878 8443
rect 1066 6789 162878 7355
rect 1066 5701 162878 6267
rect 1066 4613 162878 5179
rect 1066 3525 162878 4091
rect 1066 2437 162878 3003
<< obsli1 >>
rect 1104 2159 162840 157777
<< obsm1 >>
rect 1104 892 163286 157808
<< metal2 >>
rect 4618 0 4674 800
rect 6090 0 6146 800
rect 7562 0 7618 800
rect 9034 0 9090 800
rect 10506 0 10562 800
rect 11978 0 12034 800
rect 13450 0 13506 800
rect 14922 0 14978 800
rect 16394 0 16450 800
rect 17866 0 17922 800
rect 19338 0 19394 800
rect 20810 0 20866 800
rect 22282 0 22338 800
rect 23754 0 23810 800
rect 25226 0 25282 800
rect 26698 0 26754 800
rect 28170 0 28226 800
rect 29642 0 29698 800
rect 31114 0 31170 800
rect 32586 0 32642 800
rect 34058 0 34114 800
rect 35530 0 35586 800
rect 37002 0 37058 800
rect 38474 0 38530 800
rect 39946 0 40002 800
rect 41418 0 41474 800
rect 42890 0 42946 800
rect 44362 0 44418 800
rect 45834 0 45890 800
rect 47306 0 47362 800
rect 48778 0 48834 800
rect 50250 0 50306 800
rect 51722 0 51778 800
rect 53194 0 53250 800
rect 54666 0 54722 800
rect 56138 0 56194 800
rect 57610 0 57666 800
rect 59082 0 59138 800
rect 60554 0 60610 800
rect 62026 0 62082 800
rect 63498 0 63554 800
rect 64970 0 65026 800
rect 66442 0 66498 800
rect 67914 0 67970 800
rect 69386 0 69442 800
rect 70858 0 70914 800
rect 72330 0 72386 800
rect 73802 0 73858 800
rect 75274 0 75330 800
rect 76746 0 76802 800
rect 78218 0 78274 800
rect 79690 0 79746 800
rect 81162 0 81218 800
rect 82634 0 82690 800
rect 84106 0 84162 800
rect 85578 0 85634 800
rect 87050 0 87106 800
rect 88522 0 88578 800
rect 89994 0 90050 800
rect 91466 0 91522 800
rect 92938 0 92994 800
rect 94410 0 94466 800
rect 95882 0 95938 800
rect 97354 0 97410 800
rect 98826 0 98882 800
rect 100298 0 100354 800
rect 101770 0 101826 800
rect 103242 0 103298 800
rect 104714 0 104770 800
rect 106186 0 106242 800
rect 107658 0 107714 800
rect 109130 0 109186 800
rect 110602 0 110658 800
rect 112074 0 112130 800
rect 113546 0 113602 800
rect 115018 0 115074 800
rect 116490 0 116546 800
rect 117962 0 118018 800
rect 119434 0 119490 800
rect 120906 0 120962 800
rect 122378 0 122434 800
rect 123850 0 123906 800
rect 125322 0 125378 800
rect 126794 0 126850 800
rect 128266 0 128322 800
rect 129738 0 129794 800
rect 131210 0 131266 800
rect 132682 0 132738 800
rect 134154 0 134210 800
rect 135626 0 135682 800
rect 137098 0 137154 800
rect 138570 0 138626 800
rect 140042 0 140098 800
rect 141514 0 141570 800
rect 142986 0 143042 800
rect 144458 0 144514 800
rect 145930 0 145986 800
rect 147402 0 147458 800
rect 148874 0 148930 800
rect 150346 0 150402 800
rect 151818 0 151874 800
rect 153290 0 153346 800
rect 154762 0 154818 800
rect 156234 0 156290 800
rect 157706 0 157762 800
rect 159178 0 159234 800
<< obsm2 >>
rect 1400 856 163280 157797
rect 1400 734 4562 856
rect 4730 734 6034 856
rect 6202 734 7506 856
rect 7674 734 8978 856
rect 9146 734 10450 856
rect 10618 734 11922 856
rect 12090 734 13394 856
rect 13562 734 14866 856
rect 15034 734 16338 856
rect 16506 734 17810 856
rect 17978 734 19282 856
rect 19450 734 20754 856
rect 20922 734 22226 856
rect 22394 734 23698 856
rect 23866 734 25170 856
rect 25338 734 26642 856
rect 26810 734 28114 856
rect 28282 734 29586 856
rect 29754 734 31058 856
rect 31226 734 32530 856
rect 32698 734 34002 856
rect 34170 734 35474 856
rect 35642 734 36946 856
rect 37114 734 38418 856
rect 38586 734 39890 856
rect 40058 734 41362 856
rect 41530 734 42834 856
rect 43002 734 44306 856
rect 44474 734 45778 856
rect 45946 734 47250 856
rect 47418 734 48722 856
rect 48890 734 50194 856
rect 50362 734 51666 856
rect 51834 734 53138 856
rect 53306 734 54610 856
rect 54778 734 56082 856
rect 56250 734 57554 856
rect 57722 734 59026 856
rect 59194 734 60498 856
rect 60666 734 61970 856
rect 62138 734 63442 856
rect 63610 734 64914 856
rect 65082 734 66386 856
rect 66554 734 67858 856
rect 68026 734 69330 856
rect 69498 734 70802 856
rect 70970 734 72274 856
rect 72442 734 73746 856
rect 73914 734 75218 856
rect 75386 734 76690 856
rect 76858 734 78162 856
rect 78330 734 79634 856
rect 79802 734 81106 856
rect 81274 734 82578 856
rect 82746 734 84050 856
rect 84218 734 85522 856
rect 85690 734 86994 856
rect 87162 734 88466 856
rect 88634 734 89938 856
rect 90106 734 91410 856
rect 91578 734 92882 856
rect 93050 734 94354 856
rect 94522 734 95826 856
rect 95994 734 97298 856
rect 97466 734 98770 856
rect 98938 734 100242 856
rect 100410 734 101714 856
rect 101882 734 103186 856
rect 103354 734 104658 856
rect 104826 734 106130 856
rect 106298 734 107602 856
rect 107770 734 109074 856
rect 109242 734 110546 856
rect 110714 734 112018 856
rect 112186 734 113490 856
rect 113658 734 114962 856
rect 115130 734 116434 856
rect 116602 734 117906 856
rect 118074 734 119378 856
rect 119546 734 120850 856
rect 121018 734 122322 856
rect 122490 734 123794 856
rect 123962 734 125266 856
rect 125434 734 126738 856
rect 126906 734 128210 856
rect 128378 734 129682 856
rect 129850 734 131154 856
rect 131322 734 132626 856
rect 132794 734 134098 856
rect 134266 734 135570 856
rect 135738 734 137042 856
rect 137210 734 138514 856
rect 138682 734 139986 856
rect 140154 734 141458 856
rect 141626 734 142930 856
rect 143098 734 144402 856
rect 144570 734 145874 856
rect 146042 734 147346 856
rect 147514 734 148818 856
rect 148986 734 150290 856
rect 150458 734 151762 856
rect 151930 734 153234 856
rect 153402 734 154706 856
rect 154874 734 156178 856
rect 156346 734 157650 856
rect 157818 734 159122 856
rect 159290 734 163280 856
<< obsm3 >>
rect 3509 1123 163195 157793
<< metal4 >>
rect 4048 2128 4688 157808
rect 12208 2128 12848 157808
rect 20368 2128 21008 157808
rect 28528 2128 29168 157808
rect 36688 2128 37328 157808
rect 44848 2128 45488 157808
rect 53008 2128 53648 157808
rect 61168 2128 61808 157808
rect 69328 2128 69968 157808
rect 77488 2128 78128 157808
rect 85648 2128 86288 157808
rect 93808 2128 94448 157808
rect 101968 2128 102608 157808
rect 110128 2128 110768 157808
rect 118288 2128 118928 157808
rect 126448 2128 127088 157808
rect 134608 2128 135248 157808
rect 142768 2128 143408 157808
rect 150928 2128 151568 157808
rect 159088 2128 159728 157808
<< obsm4 >>
rect 5027 2048 12128 148749
rect 12928 2048 20288 148749
rect 21088 2048 28448 148749
rect 29248 2048 36608 148749
rect 37408 2048 44768 148749
rect 45568 2048 52928 148749
rect 53728 2048 61088 148749
rect 61888 2048 69248 148749
rect 70048 2048 77408 148749
rect 78208 2048 85568 148749
rect 86368 2048 93728 148749
rect 94528 2048 101888 148749
rect 102688 2048 110048 148749
rect 110848 2048 118208 148749
rect 119008 2048 126368 148749
rect 127168 2048 134528 148749
rect 135328 2048 142688 148749
rect 143488 2048 150848 148749
rect 151648 2048 159008 148749
rect 159808 2048 161309 148749
rect 5027 1123 161309 2048
<< labels >>
rlabel metal4 s 159088 2128 159728 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 142768 2128 143408 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 126448 2128 127088 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 110128 2128 110768 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 93808 2128 94448 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 77488 2128 78128 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 61168 2128 61808 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 44848 2128 45488 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 28528 2128 29168 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 12208 2128 12848 157808 6 VGND
port 1 nsew ground default
rlabel metal4 s 150928 2128 151568 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 134608 2128 135248 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 118288 2128 118928 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 101968 2128 102608 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 85648 2128 86288 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 69328 2128 69968 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 53008 2128 53648 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 36688 2128 37328 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 20368 2128 21008 157808 6 VPWR
port 2 nsew power default
rlabel metal4 s 4048 2128 4688 157808 6 VPWR
port 2 nsew power default
rlabel metal2 s 4618 0 4674 800 6 wb_clk_i
port 3 nsew
rlabel metal2 s 6090 0 6146 800 6 wb_rst_i
port 4 nsew
rlabel metal2 s 7562 0 7618 800 6 wbs_ack_o
port 5 nsew
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[0]
port 6 nsew
rlabel metal2 s 63498 0 63554 800 6 wbs_adr_i[10]
port 7 nsew
rlabel metal2 s 67914 0 67970 800 6 wbs_adr_i[11]
port 8 nsew
rlabel metal2 s 72330 0 72386 800 6 wbs_adr_i[12]
port 9 nsew
rlabel metal2 s 76746 0 76802 800 6 wbs_adr_i[13]
port 10 nsew
rlabel metal2 s 81162 0 81218 800 6 wbs_adr_i[14]
port 11 nsew
rlabel metal2 s 85578 0 85634 800 6 wbs_adr_i[15]
port 12 nsew
rlabel metal2 s 89994 0 90050 800 6 wbs_adr_i[16]
port 13 nsew
rlabel metal2 s 94410 0 94466 800 6 wbs_adr_i[17]
port 14 nsew
rlabel metal2 s 98826 0 98882 800 6 wbs_adr_i[18]
port 15 nsew
rlabel metal2 s 103242 0 103298 800 6 wbs_adr_i[19]
port 16 nsew
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[1]
port 17 nsew
rlabel metal2 s 107658 0 107714 800 6 wbs_adr_i[20]
port 18 nsew
rlabel metal2 s 112074 0 112130 800 6 wbs_adr_i[21]
port 19 nsew
rlabel metal2 s 116490 0 116546 800 6 wbs_adr_i[22]
port 20 nsew
rlabel metal2 s 120906 0 120962 800 6 wbs_adr_i[23]
port 21 nsew
rlabel metal2 s 125322 0 125378 800 6 wbs_adr_i[24]
port 22 nsew
rlabel metal2 s 129738 0 129794 800 6 wbs_adr_i[25]
port 23 nsew
rlabel metal2 s 134154 0 134210 800 6 wbs_adr_i[26]
port 24 nsew
rlabel metal2 s 138570 0 138626 800 6 wbs_adr_i[27]
port 25 nsew
rlabel metal2 s 142986 0 143042 800 6 wbs_adr_i[28]
port 26 nsew
rlabel metal2 s 147402 0 147458 800 6 wbs_adr_i[29]
port 27 nsew
rlabel metal2 s 25226 0 25282 800 6 wbs_adr_i[2]
port 28 nsew
rlabel metal2 s 151818 0 151874 800 6 wbs_adr_i[30]
port 29 nsew
rlabel metal2 s 156234 0 156290 800 6 wbs_adr_i[31]
port 30 nsew
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[3]
port 31 nsew
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[4]
port 32 nsew
rlabel metal2 s 41418 0 41474 800 6 wbs_adr_i[5]
port 33 nsew
rlabel metal2 s 45834 0 45890 800 6 wbs_adr_i[6]
port 34 nsew
rlabel metal2 s 50250 0 50306 800 6 wbs_adr_i[7]
port 35 nsew
rlabel metal2 s 54666 0 54722 800 6 wbs_adr_i[8]
port 36 nsew
rlabel metal2 s 59082 0 59138 800 6 wbs_adr_i[9]
port 37 nsew
rlabel metal2 s 9034 0 9090 800 6 wbs_cyc_i
port 38 nsew
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[0]
port 39 nsew
rlabel metal2 s 64970 0 65026 800 6 wbs_dat_i[10]
port 40 nsew
rlabel metal2 s 69386 0 69442 800 6 wbs_dat_i[11]
port 41 nsew
rlabel metal2 s 73802 0 73858 800 6 wbs_dat_i[12]
port 42 nsew
rlabel metal2 s 78218 0 78274 800 6 wbs_dat_i[13]
port 43 nsew
rlabel metal2 s 82634 0 82690 800 6 wbs_dat_i[14]
port 44 nsew
rlabel metal2 s 87050 0 87106 800 6 wbs_dat_i[15]
port 45 nsew
rlabel metal2 s 91466 0 91522 800 6 wbs_dat_i[16]
port 46 nsew
rlabel metal2 s 95882 0 95938 800 6 wbs_dat_i[17]
port 47 nsew
rlabel metal2 s 100298 0 100354 800 6 wbs_dat_i[18]
port 48 nsew
rlabel metal2 s 104714 0 104770 800 6 wbs_dat_i[19]
port 49 nsew
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_i[1]
port 50 nsew
rlabel metal2 s 109130 0 109186 800 6 wbs_dat_i[20]
port 51 nsew
rlabel metal2 s 113546 0 113602 800 6 wbs_dat_i[21]
port 52 nsew
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_i[22]
port 53 nsew
rlabel metal2 s 122378 0 122434 800 6 wbs_dat_i[23]
port 54 nsew
rlabel metal2 s 126794 0 126850 800 6 wbs_dat_i[24]
port 55 nsew
rlabel metal2 s 131210 0 131266 800 6 wbs_dat_i[25]
port 56 nsew
rlabel metal2 s 135626 0 135682 800 6 wbs_dat_i[26]
port 57 nsew
rlabel metal2 s 140042 0 140098 800 6 wbs_dat_i[27]
port 58 nsew
rlabel metal2 s 144458 0 144514 800 6 wbs_dat_i[28]
port 59 nsew
rlabel metal2 s 148874 0 148930 800 6 wbs_dat_i[29]
port 60 nsew
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[2]
port 61 nsew
rlabel metal2 s 153290 0 153346 800 6 wbs_dat_i[30]
port 62 nsew
rlabel metal2 s 157706 0 157762 800 6 wbs_dat_i[31]
port 63 nsew
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_i[3]
port 64 nsew
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_i[4]
port 65 nsew
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_i[5]
port 66 nsew
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_i[6]
port 67 nsew
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_i[7]
port 68 nsew
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_i[8]
port 69 nsew
rlabel metal2 s 60554 0 60610 800 6 wbs_dat_i[9]
port 70 nsew
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[0]
port 71 nsew
rlabel metal2 s 66442 0 66498 800 6 wbs_dat_o[10]
port 72 nsew
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_o[11]
port 73 nsew
rlabel metal2 s 75274 0 75330 800 6 wbs_dat_o[12]
port 74 nsew
rlabel metal2 s 79690 0 79746 800 6 wbs_dat_o[13]
port 75 nsew
rlabel metal2 s 84106 0 84162 800 6 wbs_dat_o[14]
port 76 nsew
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_o[15]
port 77 nsew
rlabel metal2 s 92938 0 92994 800 6 wbs_dat_o[16]
port 78 nsew
rlabel metal2 s 97354 0 97410 800 6 wbs_dat_o[17]
port 79 nsew
rlabel metal2 s 101770 0 101826 800 6 wbs_dat_o[18]
port 80 nsew
rlabel metal2 s 106186 0 106242 800 6 wbs_dat_o[19]
port 81 nsew
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[1]
port 82 nsew
rlabel metal2 s 110602 0 110658 800 6 wbs_dat_o[20]
port 83 nsew
rlabel metal2 s 115018 0 115074 800 6 wbs_dat_o[21]
port 84 nsew
rlabel metal2 s 119434 0 119490 800 6 wbs_dat_o[22]
port 85 nsew
rlabel metal2 s 123850 0 123906 800 6 wbs_dat_o[23]
port 86 nsew
rlabel metal2 s 128266 0 128322 800 6 wbs_dat_o[24]
port 87 nsew
rlabel metal2 s 132682 0 132738 800 6 wbs_dat_o[25]
port 88 nsew
rlabel metal2 s 137098 0 137154 800 6 wbs_dat_o[26]
port 89 nsew
rlabel metal2 s 141514 0 141570 800 6 wbs_dat_o[27]
port 90 nsew
rlabel metal2 s 145930 0 145986 800 6 wbs_dat_o[28]
port 91 nsew
rlabel metal2 s 150346 0 150402 800 6 wbs_dat_o[29]
port 92 nsew
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[2]
port 93 nsew
rlabel metal2 s 154762 0 154818 800 6 wbs_dat_o[30]
port 94 nsew
rlabel metal2 s 159178 0 159234 800 6 wbs_dat_o[31]
port 95 nsew
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[3]
port 96 nsew
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_o[4]
port 97 nsew
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[5]
port 98 nsew
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_o[6]
port 99 nsew
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_o[7]
port 100 nsew
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_o[8]
port 101 nsew
rlabel metal2 s 62026 0 62082 800 6 wbs_dat_o[9]
port 102 nsew
rlabel metal2 s 17866 0 17922 800 6 wbs_sel_i[0]
port 103 nsew
rlabel metal2 s 23754 0 23810 800 6 wbs_sel_i[1]
port 104 nsew
rlabel metal2 s 29642 0 29698 800 6 wbs_sel_i[2]
port 105 nsew
rlabel metal2 s 35530 0 35586 800 6 wbs_sel_i[3]
port 106 nsew
rlabel metal2 s 10506 0 10562 800 6 wbs_stb_i
port 107 nsew
rlabel metal2 s 11978 0 12034 800 6 wbs_we_i
port 108 nsew
<< properties >>
string FIXED_BBOX 0 0 164000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 81736714
string GDS_FILE /home/hosni/AES/caravel_aes_example/openlane/aes_example/runs/23_06_07_06_18/results/signoff/aes_example.magic.gds
string GDS_START 1593368
<< end >>

